43 years old | 0
female | 0
behavioral abnormalities (dysphoria, irritability, depressed mood) | -314,592
difficulty gaining weight | -314,592
sleep disorders (insomnia) | -314,592
increased prolactin levels | -314,592
episodes of bradycardia | -314,592
episodes of hypotension | -314,592
episodes of hypoglycemia | -314,592
cognitive problems | -314,592
poor concentration | -314,592
confusion | -314,592
memory impairment | -314,592
anxiety | -314,592
poor judgment | -314,592
carbolithium treatment | -314,592
acute onset of permanent dystonic posture | -2,184
numbness | -2,184
tingling | -2,184
diplopia | -2,184
low potassium levels | -2,184
admitted to neurology unit | -2,184
muscle relaxants treatment | -2,184
potassium treatment | -2,184
neurological bladder | -2,160
catheterized | -2,160
dystonic posture persisted | -2,160
discharged | -2,160
psychosis worsening | -2,160
carbolithium switched to olanzapine | -2,160
difficulty walking | -1,680
confined to bed | -1,680
sacral decubitus | -1,680
fever | -1,680
increased difficulty in movements | -1,680
low potassium levels | -1,680
admitted to neurology unit | -1,680
marked bradycardia | -1,680
atrial fibrillation episodes | -1,680
ventricular fibrillation episodes | -1,680
loss of consciousness | -1,680
orotracheal intubation | -1,680
transferred to intensive care unit | -1,680
involuntary parossistic eye movements | 0
involuntary head movements | 0
bilateral ptosis | 0
oculogyric crises | 0
dystonia of the head | 0
generalized muscle hypotrophy | 0
absent deep tendon reflexes | 0
normal hemocromocytometric test | 0
normal biochemical parameters | 0
normal urine analysis | 0
EEG showing diffuse theta mixed to paroxysmal activities | 0
brain MRI showing symmetric hyperintense lesions with restricted diffusion in globus pallidus | 0
episodes of bradycardia | 0
fever | 0
white blood count within 12,000 cells/μL | 0
pancytopenia | 0
procalcitonin increase (1.2 to 6.4 ng/mL) | 0
hemocultures positive for Enterococcus faecalis | 0
hemocultures positive for Acinetobacter baumanii | 0
antibiotics tigecycline infusion | 0
antibiotics colistin infusion | 0
marked bradycardia alternating with atrial fibrillation | 0
sedation required | 0
whole exome sequencing performed | 0
DDC gene mutation p.Ser250Phe (c.749C > T, rs137853208) in heterozygous state | 0
diagnosis of AADCD | 0
prescribed pyridoxine (200 mg/d) | 0
prescribed Pramipexole (0.005 mg/kg/d) | 0
sudden death | 24
abundant milk secretion after death | 24
autopsy showing sepsis | 24
no macro- and microscopic brain abnormalities | 24
