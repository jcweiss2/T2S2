73 years old | 0
male | 0
smoking | -8760
alcoholism | -8760
diabetes mellitus | -168
hypertension | -168
allergy to paracetamol | -168
no family history of hypertension | 0
no family history of diabetes mellitus | 0
no known genetic history | 0
no previous surgeries | 0
moderate to severe respiratory distress | -168
fever | -168
general malaise | -168
SARS CoV-2 positive | -168
oxygen therapy | -168
steroids | -168
no anticoagulation | -168
severe abdominal pain | -7
nausea | -7
fecal emesis | -7
fever of 39.5 °C | -7
peritoneal irritation | -7
abdominal X-ray | -7
dilated intestinal loops | -7
intestinal inter-loop edema | -7
intestinal pneumatosis | -7
admitted to hospital | 0
poor general condition | 0
frank acute abdomen | 0
radiographic data | 0
hemoglobin 15 g/dl | 0
leukocytes 17 thousand/cm3 | 0
platelets 120 thousand/cm3 | 0
procalcitonin 26 ng/ml | 0
D-dimer >5000 ng/ml | 0
high suspicion of intestinal ischemia | 0
laparotomy | 0
resection of small intestine | 0
end to end anastomosis | 0
purulent collection drained | 0
placement of drains | 0
antibiotics | 0
analgesic | 0
enoxaparin | 0
mechanical ventilation | 0
atrial fibrillation | 120
amiodarone | 120
intestinal fistula | 240
conservative treatment | 240
parenteral nutrition | 240
intestinal fistula closure | 504
pathology report | 120
ischemia and necrosis of intestinal mucosa | 120
deterioration in lung function | 720
multi-organ failure | 720
death | 720