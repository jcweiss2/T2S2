88 years old | 0
men | 0
admitted to emergency room | 0
right hemiparesis | 0
aphasia | 0
mild drowsy | 0
not communicated | 0
right hemiparesis of grade IV | 0
gaze deviation not detected | 0
visual field defect not detected | 0
diffusion-weighted MRI showed multiple small cortical infarcts | 0
atrial fibrillation | -5184
hypertension | -5184
hyperlipidemia | -5184
gout | -5184
chronic renal insufficiency | -5184
old basal ganglia lacunar infarct | -5184
antiplatelet agent | -5184
medication for permanent atrial fibrillation not administered | -5184
multiple small cortical infarcts in left middle cerebral artery territory | 0
involvement of insular cortex not detected | 0
electrocardiogram revealed atrial fibrillation with rapid ventricular rhythm | 0
echocardiogram revealed moderate aortic valve regurgitation | 0
left atrial enlargement | 0
ejection fraction normal | 0
thrombus not observed in the atrium or ventricle | 0
treatment with heparin | 0
treatment with digoxin | 0
digoxin stopped | 48
anticoagulation stopped | 168
gross hematuria | 168
intubation performed | 432
purulent sputum | 432
severe stridor | 432
epiglottitis | 432
right-sided weakness progressed to hemiplegia | 432
consciousness decreased to stuporous state | 720
eyeball deviated to right side | 720
left side hemiparesis of grade I | 720
diffuse subcortical infarcts of middle cerebral artery territory | 720
insular cortex not directly involved | 720
atrial fibrillation converted to normal sinus rhythm | 720
cardiac enzymes normal | 720
follow-up echocardiogram not different | 720
normal sinus rhythm sustained | 720
died due to sepsis | 831
second ischemic attack | 720
first attack | 0 
second cerebral infarct | 720 
first cerebral infarct | 0 
sepsis | 831