62 years old | 0
female | 0
headache | -96
fever | -96
rigor | -96
Pfizer COVID-19 vaccine | -120
ceftriaxone allergy | 0
disorientation | 0
inability to talk | 0
meningeal irritation signs | 0
isocor pupils | 0
positive light reaction | 0
Babinski sign | 0
inability to stand | 0
inability to walk | 0
wheelchair use |> 0
elevated body temperature | 0
temp. 38C | 0
SPO2 98% | 0
pulse rate 105 bpm | 0
blood pressure 125/80 mmHg | 0
mild leukocytosis | 0
agranulocytosis | 0
elevated CRP | 0
normal serum electrolyte | 0
normal renal function tests | 0
normal liver function tests | 0
random blood sugar 185mg/dl | 0
normal brain CT scan | 0
normal brain MRI | 12
clear CSF | 12
lymphocytic pleocytosis | 12
protein 802mg/dl | 12
glucose 71mg/dl | 12
lactate 19.61mg/dl | 12
negative gram stain | 12
negative Herpes simplex PCR | 12
meropenem IV | -96
dexamethasone IV | -96
acyclovir IV | 0
consciousness restored | 48
oriented | 48
discharged | 336
