74 years old | 0
woman | 0
newly diagnosed diabetes mellitus | -504
hypertension | -?
hyperlipidemia | -?
small cell lung cancer metastatic to the brain | -504
presented to the emergency department | 0
lethargy | -48
weakness | -48
significantly worsened over the past 2 days | -48
cancer diagnosed | -504
gamma knife radiation therapy | -504
dexamethasone 4 mg twice daily | -504
cerebral edema | -504
diabetes mellitus diagnosed | -504
hemoglobin A1c 6.5% | -504
blood glucose >799 mg/dL | 0
hemoglobin A1c 10.8% | 0
follow-up appointment with oncologist | -?
blood glucose elevated | -?
no symptoms | -?
advised to follow up with primary care provider | -?
started to feel ill | -?
went to ED instead | 0
admitted with hyperosmolar hyperglycemic state | 0
left eyelid swelling | 0
erythema | 0
preseptal cellulitis | 0
ophthalmoplegia | 0
visual impairment left eye | 0
worsened mental status | 0
difficulty following commands | 0
aggressive hydration with IV fluids | 0
insulin | 0
septic shock | 0
broad-spectrum antibiotics | 0
vasopressors via central venous catheter | 0
evaluated in medical ICU | ?
poor prognosis | 0
not a candidate for ICU-level care | 0
medically managed on inpatient medicine service | 0
computed tomography scan head and neck | 0
left ocular proptosis | 0
invasive rhinomaxillary fungal disease | 0
amphotericin B started | 0
urgent surgical debridement | 0
magnetic resonance imaging head and neck | ?
invasive fungal disease left inferior frontal lobe | 0
multidisciplinary meeting | ?
healthcare agent declined further surgery | ?
orbital exenteration offered | ?
skull base surgery offered | ?
healthcare agent preferred conservative medical management | ?
surgical pathology confirmed invasive mucormycosis (R. oryzae) | ?
concomitant infection S. maltophilia | ?
blood cultures grew methicillin-susceptible S. aureus | ?
treated with liposomal amphotericin B | 0
cefazolin | 0
levofloxacin | 0
herpetic lesion | ?
resolved with valacyclovir | ?
vasopressor support until hospital day 19 | 19 * 24 = 456
electrolyte abnormalities | 0
hypokalemia | 0
pronounced after liposomal amphotericin B started on day 5 | 5 * 24 = 120
potassium level 4.2 mmol/L | 0
hypokalemia persisted | 120
potassium supplementation | 120
spironolactone | 120
completed course on day 25 | 25 * 24 = 600
discharged day 26 | 26 * 24 = 624
lost to follow-up | 624
declined appointments | 624
hypertension | -504
hyperlipidemia | -504
gamma knife radiation therapy | -336
dexamethasone 4 mg twice daily | -336
cerebral edema | -336
follow-up appointment with oncologist | -120
blood glucose elevated | -120
no symptoms | -120
advised to follow up with primary care provider | -120
started to feel ill | -24
difficulty following commands |> 0
evaluated in medical ICU | 96
poor prognosis | 96
not a candidate for ICU-level care | 96
amphotericin B started | 120
urgent surgical debridement | 120
magnetic resonance imaging head and neck | 120
invasive fungal disease left inferior frontal lobe | 120
multidisciplinary meeting | 120
healthcare agent declined further surgery | 120
orbital exenteration offered | 120
