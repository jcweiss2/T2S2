20 years old | 0
African American | 0
female | 0
weight 75 kg | 0
height 1.75 meters | 0
body mass index 24.5 kg.m-2 | 0
admitted | 0
postictal state | 0
generalized tonic-clonic seizure | 0
new-onset headache | 0
blood pressures 170–140 mmHg | 0
blood pressures 120–90 mmHg | 0
prenatal care unremarkable | 0
medical history negative for hypertensive disorders | 0
medical history negative for seizure disorders | 0
platelet count 124,000 per cubic millimeter | 0
alkaline phosphatase 207 IU.L-1 | 0
alanine aminotransferase 60 IU.L-1 | 0
aspartate aminotransferase 50 IU.L-1 | 0
lactate dehydrogenase 353 IU.L%1 | 0
uric acid 7.4 mg.dL-1 | 0
Prothrombin Time 9.9 seconds | 0
fibrinogen 463 mg.dL-1 | 0
3+ urine protein | 0
International Normalized Ratio 0.9 | 0
Partial Thromboplastin Time 29.2 seconds | 0
magnesium sulfate infusion started | 0
neurological checks | 0
blood tests | 0
continuous fetal monitoring | 0
clinical stabilization | 0
blood pressures 160–140 mmHg | 0
blood pressures 100–80 mmHg | 0
neurologically improving | 0
awake | 0
alert | 0
responsive | 0
oriented | 0
intact motor strength | 0
intact sensations | 0
no more seizure episodes | 0
denied headache | 0
denied visual disturbances | 0
betamethasone received | 0
clinically stable | 0
reassuring fetal status | 0
platelet count decreased to 97,000 per cubic millimeter | -3
HELLP syndrome possibility | -3
repeat coagulation profile | -3
low PT | -3
elevated fibrinogen | -3
normal INR | -3
normal PTT | -3
risk of recurrent seizures | -3
risk of disseminated intravascular coagulation | -3
risk of stroke | -3
cesarean section decided | -3
Thromboelastography performed | -3
Reaction time 5.8 minutes | -3
Kinetics time 1.8 minutes | -3
alpha angle 66.2 degrees | -3
Lysis index 30 (LY30) 0% | -3
Maximal Amplitude 66.2 mm | -3
spinal anesthesia performed | 0
hyperbaric 0.75% bupivacaine 14.25 mg | 0
intrathecal morphine 0.02 mg | 0
lumbar 3–4 intervertebral space | 0
adequate thoracic 4-sensory level block | 0
cesarean section uneventful | 0
neonate APGAR scores 7/7/7 | 0
neonatal intensive care unit admission | 0
hemodynamically stable | 0
blood pressures 140–130 mmHg | 0
blood pressures 90–60 mmHg | 0
magnesium infusion continued | 0
no cardiovascular supportive medications | 0
blood loss 700 mL | 0
recovery unremarkable | 0
post-spinal anesthesia evaluation unremarkable | 0
no neuraxial hematoma | 0
platelet counts improved | 24
liver function tests improved | 24
discharged | 120
