57 years old | 0
    man | 0
    brought unconscious to Emergency Department | 0
    abuse alcohol | 0
    alcohol dementia | 0
    arterial hypertension | 0
    fully conscious | -24
    increasingly confused | -12
    unresponsive | -6
    previous hospitalization after intake of antifreeze coolant | -672
    ethylene glycol poisoning suspected | -672
    ethylene glycol poisoning confirmed | -672
    Glasgow coma scale 3/15 | 0
    cyanotic | 0
    hypothermic (temperature 34.7°C) | 0
    Kussmaul breathing (28 breaths per min) | 0
    blood pressure 150/90 mmHg | 0
    heart rate fluctuating (75–150 beats per min) | 0
    atrial fibrillation (92 beats per min) | 0
    no ECG abnormalities | 0
    rigid limbs | 0
    pupils with absent light reflex | 0
    computed tomography of cerebrum unremarkable | 0
    chest X-ray unremarkable | 0
    hyperkalemia (K+=5.1 mmol/L) | 0
    high anion gap (34.7 mEq/L) | 0
    elevated lactic acid (>30 mmol/L) | 0
    arterial blood gas test: pH 7.07 | 0
    arterial blood gas test: HCO3− 6.4 mmol/L | 0
    bladder catheterization: clear urine | 0
    urine drug screening positive for benzodiazepines | 0
    intubated | 0
    transmitted to ICU | 0
    treatment with bicarbonate | 0
    electrolyte correction | 0
    intravenous ethyl alcohol infusion | 0
    suspicion of sepsis | 0
    intravenous antibiotics (Meropenem and Metronidazole) | 0
    first signs of renal failure | 6
    increasing creatinine (90 to 138 µmol/L) | 6
    decreasing urine production | 6
    hyperkalemia | 6
    worsening acidosis (pH 6.90) | 6
    increased anion gap (35.5 mEq/L) | 6
    hemodialysis initiated | 6
    hypotension | 6
    increased heart rate | 6
    urine sediment examination showing COM crystals | 6
    clinical recovery | 48
    extubated | 48
    hemodialysis discontinued | 48
    ethyl alcohol infusion discontinued | 48
    acceptable urine production under furosemide | 48
    normalized creatinine | 48
    normalized calcium | 48
    corrected acidosis | 48
    decreasing lactate | 48
    transferred to medical ward | 48
    discharged | 48
