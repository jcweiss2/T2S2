66 years old | 0  
    male | 0  
    hypertension | 0  
    hyperlipidemia | 0  
    hepatitis C virus infection | 0  
    atrial fibrillation | 0  
    anticoagulated with apixaban | 0  
    fall | 0  
    dizziness | 0  
    lost consciousness | 0  
    found down | 0  
    Glasgow Coma Score of 15 | 0  
    no focal neurological deficits | 0  
    noncontrast CT head | 0  
    right frontal subdural hematoma | 0  
    right medial orbital wall fracture | 0  
    minimal mass effect | 0  
    admitted to surgical intensive care unit | 0  
    severe headache | 24  
    head CT repeated | 24  
    worsening subdural hematoma | 24  
    associated mass effect | 24  
    2 mm midline shift | 24  
    remained neurologically intact | 24  
    discharged to acute inpatient rehabilitation | 144  
    repeat head CT in 2 weeks | 144  
    terrible headache | 168  
    repeat neurosurgical evaluation | 168  
    neurologically intact | 168  
    repeat CT head | 168  
    expansion of hematoma to 15 mm | 168  
    increased mass effect | 168  
    8 mm midline shift | 168  
    underwent burr holes for evacuation | 168  
    placement of subdural drain | 168  
    headache improved | 168  
    SDH decreased in size | 168  
    drain removed | 216  
    discharged home | 216  
    levetiracetam for seizure prophylaxis | 216  
    strange sensation in right arm | 360  
    feeling of inability to control arm | 360  
    sent to emergency room | 360  
    focal left arm seizure | 360  
    treated for seizure | 360  
    started on EEG monitoring | 360  
    admitted | 360  
    unresponsive | 384  
    CT head showed no acute hemorrhage | 384  
    EEG indicated status epilepticus | 384  
    intubated | 384  
    transferred to medical intensive care unit | 384  
    cerebral CTA obtained | 384  
    negative for pathology | 384  
    ventilator-dependent respiratory failure | 384  
    septic shock secondary to Pseudomonas bacteremia | 384  
    tracheostomy | 384  
    gastrostomy | 384  
    stabilized | 384  
    discharged to long-term acute care hospital | 696  
    levetiracetam | 696  
    oxcarbazepine | 696  
    less responsive | 744  
    transferred back for neurosurgical evaluation | 744  
    opened eyes to stimulation | 744  
    localized with right upper extremity | 744  
    minimal movement of left upper and bilateral lower extremities | 744  
    cough | 744  
    gag | 744  
    corneal reflexes | 744  
    pupillary reflexes | 744  
    CT and CTA head | 744  
    right frontal intraparenchymal hemorrhage | 744  
    no vascular lesion or anomaly | 744  
    cerebral catheter angiography performed | 744  
    prominence of anterior temporal branch of right middle cerebral artery | 744  
    early shunting of blood through cortical vein | 744  
    opacification of capillary-like serpiginous tangle of vessels | 744  
    AVM Spetzler-Martin Grade 1 | 744  
    AVM Spetzler-Ponce Grade A | 744  
    embolization of AVM performed | 768  
    embolization successful | 768  
    no opacification of draining vein | 768  
    no AVM nidus seen | 768  
    taken to operating room for resection | 912  
    right pterional craniotomy performed | 912  
    AVM separated from surrounding parenchyma | 912  
    feeding arteries coagulated | 912  
    draining vein coagulated | 912  
    resection | 912  
    intraoperative Doppler ultrasound | 912  
    no arterial flow in draining vein | 912  
    intraparenchymal hematoma evacuated | 912  
    postoperative angiography | 912  
    no residual AVM | 912  
    mental status progressively improved | 936  
    followed commands | 936  
    tracked with eyes | 936  
    spontaneous antigravity movement of right upper extremity | 936  
    no movement of left upper or bilateral lower extremities | 936  
    postoperative course complicated by Pseudomonas sepsis | 936  
    treated by infectious disease | 936  
    discharged to long-term acute care | 1080  
