26 years old | 0
female | 0
admitted to the hospital | 0
headache | -336
nonresponsive to anti-inflammatory drugs | -336
right-sided weakness | 0
visual disturbances | 0
combined (estrogen-progestogen) contraceptives | -8760
ChAdOx1 nCoV-19 vaccine | -336
severe right-sided weakness | 0
no visual field defects | 0
hyperdense rectus sinus and vein of Galen | 0
multifocal venous thrombosis | 0
bilateral occlusion of parietal cortical veins | 0
straight sinus, vein of Galen, internal cerebral veins and inferior sagittal sinus | 0
transverse sinuses partially involved | 0
extensive venous infarction with hemorrhagic transformation | 0
D-dimer dramatically raised | 0
platelet count 134x10^9/L | 0
fondaparinux | 0
decreased consciousness | 24
right-sided hemiplegia | 24
complete Balint syndrome | 24
IVIG | 24
dexamethasone | 24
argatroban | 24
neurological conditions improved | 48
right upper-limb strength recovered | 48
partial optic ataxia | 48
regression of apraxia | 48
rectus sinus and vein of Galen normal density | 144
oedema in brain tissue | 144
restored venous flow in rectus sinus and vein of Galen | 168
right internal cerebral vein and bilateral frontoparietal cortical veins still occluded | 168
large intraparenchimal venous infarction unchanged | 168
platelet count increased to 339x10^9/L | 168
D-dimer decreased to normal levels | 168
aPF4 reactivity reduced | 168
moderate disability | 1440
no neuropsychological deficits | 1440
can walk unassisted for short distances | 1440
sustained clonus and spasticity in right leg | 1440
right arm almost fully recovered | 1440
fondaparinux replaced with oral vitamin K antagonist | 1440