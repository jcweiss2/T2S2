17 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
Caucasian | 0 | 0 | Factual
throat pain | -168 | 0 | Factual
odynophagia | -168 | 0 | Factual
blood tests | -168 | -168 | Factual
Hemoglobin: 7.0 g/dL | -168 | -168 | Factual
Hematocrit: 21% | -168 | -168 | Factual
WBC: 33 x 10^9 cells/L | -168 | -168 | Factual
platelets: 38 x 10^9 cells/L | -168 | -168 | Factual
Acute promyelocytic leukemia (M3) | -168 | -168 | Factual
daunorubicin | -168 | 0 | Factual
vesanoid | -168 | 0 | Factual
necrotic lesion | 0 | 0 | Factual
unpleasant odor | 0 | 0 | Factual
biopsy | 0 | 0 | Factual
culture | 0 | 0 | Factual
nonspecific chronic diffuse inflammation | 0 | 0 | Factual
necrotic areas | 0 | 0 | Factual
numerous bacteria | 0 | 0 | Factual
Enterococcus spp | 0 | 0 | Factual
Staphylococcus aureus | 0 | 0 | Factual
Candida SP | 0 | 0 | Factual
noma-like lesion | 0 | 0 | Factual
antibiotic therapy | 0 | 45 | Factual
ceftazidime | 0 | 45 | Factual
amicacin | 0 | 45 | Factual
vancomycin | 0 | 45 | Factual
fluconazole | 0 | 45 | Factual
penicillin G | 0 | 45 | Factual
pneumonia | 0 | 45 | Factual
sepsis | 0 | 45 | Factual
intensive care unit | 0 | 45 | Factual
total recovery | 45 | 45 | Factual
extensive loss of soft palate tissue | 45 | 45 | Factual
mucocutaneous leishmaniasis | 0 | 0 | Negated
lupus erythematosus | 0 | 0 | Negated
leprosy | 0 | 0 | Negated
agranulocytic ulcerations | 0 | 0 | Negated
physical trauma | 0 | 0 | Negated
syphilis | 0 | 0 | Negated
oral cancer | 0 | 0 | Negated
yaws | 0 | 0 | Negated