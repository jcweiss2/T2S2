26 years old | 0
female | 0
laparoscopic cholecystectomy | -672
lump in right upper quadrant | 0
malaena episodes | 0
pale | 0
anicteric | 0
pulse rate 120/min | 0
blood pressure 90/60 mmHg | 0
respiratory rate 25/min | 0
tender lump in right upper quadrant | 0
progressive pallor | 8
hypotension | 8
malena episodes | 8
emergency ultrasound | 8
free fluid in lower abdomen | 8
encysted collection around liver | 8
bidirectional flow pattern on Doppler | 8
CT abdomen with vascular reconstruction | 8
hemoglobin 5.6 g/dl | 8
elevated hepatic enzymes | 8
normal coagulation profile | 8
IV fluids resuscitation | 8
packed red blood cells transfusion | 8
perihepatic collection | 8
contrast spillage in gallbladder fossa | 8
HAPA involving right hepatic artery | 8
deterioration despite resuscitation | 24
exploratory laparotomy | 24
right subcostal incision | 24
evacuation of clotted blood | 24
isolation of right hepatic artery | 24
control of proximal artery | 24
rupture of pseudoaneurysmal sac | 24
excision of pseudoaneurysmal sac | 24
identification of pseudoaneurysm in cystic artery stump | 24
metal clip erosion in right hepatic artery | 24
repair of right hepatic artery rent | 24
peritoneal lavage | 24
wide bore drain placement | 24
haemostasis | 24
wound closure in two layers | 24
post-operative packed red blood cells transfusion | 24
superficial surgical site infection | 288
wound dressings | 288
discharge | 288
no delayed biliary stricture | 2160
no liver dysfunction | 2160
bidirectional flow on ultrasound | 2160
planned follow-up for 2 years | 2160
