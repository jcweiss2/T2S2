62 years old | 0
male | 0
ankle twisting injury | -48
undisplaced fracture medial malleolus | -48
below knee ankle plaster (slab) | -48
advised elevation | -48
medical history negative for diabetes | 0
medical history negative for allergic conditions | 0
analgesic with proteolytic | -48
itching | -12
pain | -12
swelling | -12
erythema up to distal thigh | -12
slab removed | -12
fever | -12
progressive swelling | -12
crepitus | -12
blisters getting peeled off easily | -12
serous discharge | -12
sequential discoloration of tissue from pinkish to velvety | -12
blackening due to necrosis | -12
foul smell | -12
necrotizing fasciitis diagnosis | -12
referred to tertiary care center | 24
2 cm incision in the skin down to deep fascia | 96
lack of bleeding | 96
dishwater-colored fluid seeping from the wound | 96
positive finger probe test | 96
Pseudomonas aeruginosa cultured | 96
gas gangrene ruled out | 96
Pseudomonas resistant to piperazillin-tazobactam | 96
meropenem switched | 96
teicoplanin switched | 96
clindamycin switched | 96
above knee amputation | 168
necrotizing fasciitis continued to expand above stump | 168
debridement on day 9 | 216
debridement on day 12 | 288
debridement on day 15 | 360
septic shock | 480
acute renal failure | 480
death | 480
