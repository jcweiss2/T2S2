50 years old | 0
female | 0
admitted to the emergency department | 0
epigastric pain | -360
fever | -360
chill | -360
nausea | -360
abdominal surgery for multiple biliary stones | -19200
history of choledochoduodenostomy | -19200
acute, continuous, dull-like pain | 0
tender on the right upper quadrant area | 0
white blood cell count, 14,760/mm3 | 0
hemoglobin level, 10.0 g/dL | 0
erythrocyte sedimentation ratio, 140 mm/hr | 0
c-reactive protein level, 23.89 mg/dL | 0
aspartate aminotransferase level (AST), 101 IU/L | 0
alanine aminotransferase (ALT) level, 114 IU/L | 0
total billirubin, 4.6 mg/dL | 0
amylase level, 48 U/L | 0
abdominal computed tomographic (CT) scan | 0
multiple stones in the common bile duct (CBD) and intra-hepatic duct (IHD) | 0
biliary obstruction | 0
multifocal liver abscesses | 0
air-biliarygram | 0
emergency ERCP | 0
opening of a choledochoduodenostomy | 0
cholangiogram | 0
multiple filling defects in the CBD | 0
extraction of brown-pigmented mud stones | 1
hypoxic | 2
bradycardic | 2
comatose | 3
cardiac arrest | 3
termination of the procedure | 3
cardio-pulmonary resuscitation | 3
intubation | 3
transfer to the intensive care unit | 4
death | 5
massive systemic air embolism | 5
biliary-venous fistula | 5
choledochoduodenostomy | -19200 
liver abscesses | -360 
ERCP | 0 
sphincterotomy | 0 
percutaneous transhepatic biliary drainage (PTBD) | 0 
high intraluminal air pressure | 0 
air embolism | 2 
cardio-pulmonary system | 5 
fatal air embolism | 5 
liver biopsy | 0 
hepatobiliary system | 0 
barotraumas | 0 
multiple liver abscesses | 0 
insufflated air | 0 
massive air embolisms | 5 
abrupt deterioration of vital and neurologic signs | 2 
chest X-ray | 5 
air density occupied in heart chambers | 5 
hepatic vasculatures and splenic vein | 5 
air embolism in the cardio-pulmonary system | 5