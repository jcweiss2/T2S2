60 years old | 0
female | 0
admitted to the hospital | 0
right otalgia | -72
purulent otorrhea | -72
right malignant otitis externa | 0
intravenous Augmentin | 0
refractory to antibiotic treatment | 120
computed tomography scan of the right temporal bone | 120
bony destruction of external auditory canal | 120
mastoid destruction | 120
right mandibular fossa destruction | 120
osteomyelitis of the right temporal bone | 120
severe sepsis | 192
metabolic acidosis | 192
acute renal failure | 192
intubated | 192
managed in the surgical intensive care unit | 192
multi-resistant Staphylococcus aureus | 192
Pseudomonas aeruginosa | 192
Candida albicans | 192
intravenous meropenem | 192
intravenous vancomycin | 192
intravenous caspofungin | 192
anuric | 192
dialysis | 192
sustained low efficiency dialysis | 192
continuous venoE veno-venous hemodialysis | 192
abdominal distension | 264
abdominal X-ray | 264
mottled lucencies over the gastric lumen | 264
computed tomography scan of the abdomen and pelvis | 264
extensive gastric intramural gas | 264
exploratory laparotomy | 264
infarcted stomach from the cardia to the pylorus | 264
total gastrectomy | 264
palpable pulsations of coeliac axis and superior mesenteric artery | 264
persistent hypotension | 336
bradycardia | 336
maximal inotropic support | 336
passed away | 408
total gastric infarction | 264
widely disseminated fungal organisms | 264
infarction of the entire gastric wall | 264
ghost outline preservation of architectural features | 264
fungal organisms disseminated through the entire gastric wall | 264
fungal spores and hyphae | 264
branching at right angles | 264
mucormycosis | 264
arterial thrombosis | 264
tissue infarction | 264
necrosis | 264
venous invasion | 264
hemorrhage | 264
resistant to anti-fungal agents | 336
angioinvasion | 336
thrombosis of vessels | 336
less optimal penetration of medications | 336
