67 years old | 0
    male | 0
    hypertension | -876000
    benign prostatic hyperplasia | -876000
    childhood asthma | -876000
    abdominal pain | -672
    bloating | -672
    decreased oral intake | -672
    shortness of breath | -672
    fatigue | -672
    no bowel movement | -72
    no fever | 0
    no chills | 0
    no cough | 0
    no trauma | 0
    no weight loss | 0
    no nausea | 0
    no vomiting | 0
    no diarrhea | 0
    no sick contacts | 0
    no recent travel | 0
    no hematuria | 0
    no hematochezia | 0
    no new diet | 0
    no unusual foods | 0
    retired office manager | 0
    former smoker | 0
    drinking two to three beers daily | 0
    finasteride | 0
    omeprazole | 0
    tamsulosin | 0
    afebrile | 0
    blood pressure 102/47 mm Hg | 0
    heart rate 149 beats per minute | 0
    saturating well on room air | 0
    bilateral decreased breath sounds | 0
    wheezing at bases | 0
    tachycardia | 0
    irregularly irregular pulse | 0
    trace bilateral pedal edema | 0
    soft abdomen | 0
    mildly distended abdomen | 0
    diffuse tenderness | 0
    atrial fibrillation with rapid ventricular rate | 0
    elevated white blood count | 0
    ProBNP 11,442 pg/mL | 0
    negative COVID-19 test | 0
    creatinine 1.84 mg/dL | 0
    elevated D-dimer 6.45 mg/L | 0
    chest X-ray minimal infiltrates | 0
    chest X-ray cardiomegaly | 0
    chest X-ray mild pleural effusion bilaterally | 0
    echocardiogram normal ejection fraction | 0
    echocardiogram no right heart strain | 0
    CT angiography positive for right lower lobe pulmonary embolism | 0
    CT angiography mild abdominal ascites | 0
    CT abdomen extensive abdominal and pelvic ascites | 0
    CT abdomen no bowel obstruction | 0
    CT abdomen unremarkable liver morphology | 0
    prophylactic antibiotic coverage | 0
    admitted to intensive care unit | 0
    negative urine culture | 0
    negative blood culture | 0
    abdominal discomfort persisted | 0
    afib RVR managed | 0
    anticoagulated for PE | 0
    worsening abdominal distension | 0
    paracentesis completed twice | 0
    initial paracentesis 4250 cc straw-colored fluid | 0
    ascitic fluid analysis no spontaneous bacterial peritonitis | 0
    ascitic fluid pathology atypical epithelioid cells | 0
    viral hepatitis serologies noncontributory | 0
    liver function tests noncontributory | 0
    Alpha-fetoprotein noncontributory | 0
    CA 19-9 noncontributory | 0
    CEA noncontributory | 0
    ANA noncontributory | 0
    anti-smooth muscle antibody noncontributory | 0
    anti-mitochondrial antibody noncontributory | 0
    SAAG 0.8 | 0
    family history reviewed | 0
    social history reviewed | 0
    no asbestos exposure | 0
    worked in rum factory administrative capacity | 0
    new-onset nausea | 168
    new-onset vomiting | 168
    new-onset diarrhea | 168
    repeat CT abdomen/pelvis multiple dilated loops of small bowel | 168
    repeat CT abdomen/pelvis high-grade small bowel obstruction | 168
    repeat CT abdomen/pelvis thickened omentum | 168
    repeat CT abdomen/pelvis questionable peritoneal carcinomatosis | 168
    exploratory laparotomy | 168
    advanced carcinomatosis | 168
    matted visceral structures | 168
    probable malignant ascites | 168
    rapid decompensation | 360
    expired | 360
    final pathology primary MPM | 360
    abdominal fluid malignant mesothelioma | 360
    immunohistochemistry mesothelial phenotypic expression | 360
    peritoneum excision malignant epithelioid mesothelioma | 360
    rhabdoid features | 360
    