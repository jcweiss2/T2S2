76 years old|0
male|0
admitted to the emergency department for severe hyponatremia|0
medical history includes pancreatic adenocarcinoma with metastasis to the liver|0
diastolic heart failure|0
atrial fibrillation|0
coronary artery disease|0
scheduled to undergo port placement for chemotherapy|0
sodium level of 116 mmol/L|0
sent to the emergency department for further evaluation|0
x-ray findings consistent with pneumonia|0
started on broad-spectrum antibiotics|0
receiving small boluses of fluid for hyponatremia|0
transferred to the intensive care unit|0
jugular vein distention|0
lower extremity pitting edema|0
transthoracic echocardiogram (TTE) ordered|0
normal left ventricular cavity size|0
mildly reduced systolic function|0
septal flattening|0
left atrial enlargement|0
suspected MV vegetation|0
severe mitral regurgitation|0
tricuspid regurgitation Doppler confirmed an elevated RV systolic pressure|0
elevated right heart pressure attributed to type 2 and type 3 pulmonary arterial hypertension|0
ill-defined thickening in the TV leaflets|0
afebrile|0
leukocytosis|0
history of recent urethral instrumentation for a urological procedure|0
blood cultures obtained on day 1|0
infectious disease specialist consulted|0
continued on broad-spectrum antibiotics|0
scheduled for a transesophageal echocardiogram (TEE) the following day|0
TEE showed normal left ventricular size and function|24
ejection fraction of 60%-65%|24
normal RV size and function|24
hypermobile interatrial septum without patent foramen ovale|24
no left atrial or left atrial appendage thrombus|24
2 large vegetations on the atrial aspect of MV leaflets|24
anterior leaflet measuring 1.3 × 1.1 cm|24
posterior leaflet measuring 1.2 × 0.9 cm|24
severe mitral regurgitation with systolic flow reversal in the pulmonary vein|24
large 1.6 × 1.1 cm vegetation on the TV leaflet|24
tricuspid regurgitation|24
RVSP 47 mm Hg|24
blood cultures negative for growth on 4 repeat cultures|24
polymerase chain reaction testing for Coxiella urnetiid, Legionella spp, and Brucella spp negative|24
workup for antiphospholipid syndrome unremarkable|24
presence of vegetations on both the MV and TV|24
persistently negative blood cultures|24
metastatic pancreatic cancer|24
suspected diagnosis of marantic endocarditis|24
previously treated with apixaban|0
apixaban discontinued due to severe thrombocytopenia|24
recommended to start on low molecular weight heparin or unfractionated heparin|24
computed tomography imaging of the head completed|24
discontinued from broad-spectrum antibiotics|24
observation of clinic course to clarify diagnosis|24
started on enoxaparin once platelets recovered above 50,000 109/L|24
patient expired shortly after discovery of valvular regurgitation|24
death within weeks of discharge|24
