28 years old | 0
    woman | 0
    hypochondriac pain | -840
    pain radiating to the back | -840
    jaundice | -672
    tea-colored urine | -672
    no known medical illness | 0
    no history of surgery | 0
    blood pressure 145/94 mm Hg | 0
    pulse rate 80 bpm | 0
    afebrile | 0
    hyperbilirubinaemia | 0
    ALT normal | 0
    AST normal | 0
    ALP normal | 0
    white cell count 8.6×10^9/L | 0
    normal renal profile | 0
    normal coagulation profile | 0
    normal serum amylase | 0
    gallstone | 0
    no dilated biliary ducts | 0
    bilirubin increased from 57.6 μmol/L to 126.4 μmol/L | 0
    ALP increased from 237 units/L to 357 units/L | 0
    ALT increased from 251 units/L to 523 units/L | 0
    AST increased from 266 units/L to 288 units/L | 0
    no fever | 0
    dilated intrahepatic biliary ducts | 0
    dilated extrahepatic biliary ducts | 0
    lesion in the distal bile duct | 0
    diagnosis of impacted soft stone in the common bile duct | 0
    referred for emergency ERCP | 0
    denied travel | 0
    denied contact with COVID-19 positive individuals | 0
    denied COVID-19 symptoms | 0
    signed health declaration | 0
    not tested for COVID-19 | 0
    staff screened for COVID-19 | 0
    health declaration by staff | 0
    protocol checklist for endoscopy | 0
    patient arrival to institution | 0
    body temperature check | 0
    staff wearing surgical masks | 0
    hand hygiene | 0
    patient sent to operating theatre | 0
    patient wearing waterproof gown | 0
    checklist for conscious sedation | 0
    intravenous antibiotic administered | 0
    seven staff involved in ERCP | 0
    radiation precautions | 0
    donning PPE | 0
    hand hygiene before donning | 0
    N95 respirator | 0
    visor | 0
    lead shield aprons | 0
    thyroid shields | 0
    disposable OT gown | 0
    double gloves | 0
    patient positioned prone | 0
    oxygen therapy | 0
    vital signs monitored | 0
    intravenous sedative | 0
    protective barrier applied | 0
    transparent plastic sheet for communication | 0
    scope entry slit | 0
    Yankauer sucker slit | 0
    ampulla floppy | 0
    pus observed | 0
    partial sphincterotomy | 0
    guide wire in bile duct | 0
    10-French stent deployed | 0
    bile flow good | 0
    reversal medication administered | 0
    patient awake | 0
    endoscopy equipment disinfection | 0
    doffing PPE | 0
    removal of gloves | 0
    gown removal | 0
    visor disinfection | 0
    mask removal | 0
    new mask applied | 0
    shoe cover removal | 0
    hand hygiene post-doffing | 0
    patient cleaning | 0
    gown removal | 0
    cap change | 0
    new mask applied | 0
    patient transferred to recovery | 0
    intravenous antibiotics continued | 0
    equipment disinfection | 0
    floor disinfection | 0
    surface disinfection | 0
    bilirubin decreased to 50 μmol/L | 72
    leucocyte count 9.98×10^9/L | 72
    ALP decreased to 354 units/L | 72
    ALT decreased to 359 units/L | 72
    AST decreased to 100 units/L | 72
    discharged after 5 days | 120
    bilirubin 21.8 μmol/L | 336
    ALP 134 units/L | 336
    ALT 21 units/L | 336
    AST 20 units/L | 336
    scheduled for ERCP in 6 weeks | 336

    