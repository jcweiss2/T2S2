62 years old | 0
    man | 0
    brought to the emergency department | 0
    found unresponsive in bed | 0
    wife reported 5-day history of bilateral otalgia | -120
    not improved by use of olive oil ear drops | -120
    presumed impacted ear wax | -120
    Glasgow Coma Scale score at scene was 8 | -120
    past medical history included CRS with nasal polyposis | -120
    previously underwent functional endoscopic sinus surgery | -120
    nasal polypectomy | -120
    chronic obstructive pulmonary disease | -120
    hypertension | -120
    glaucoma | -120
    right sided keratoconus treated with previous corneal graft | -120
    hypercholesterolaemia | -120
    regular medications included beclomethasone/formoterol inhaler | -120
    salbutamol inhaler | -120
    amlodipine | -120
    simvastatin | -120
    beclometasone dipropionate nasal spray | -120
    examination: tachypnoeic (25 breaths per minute) | 0
    tachycardic (120 beats per minute) | 0
    pyrexial (40°C) | 0
    Glasgow Coma Scale was 11 | 0
    bilateral green purulent rhinorrhea | 0
    bilateral proptosis | 0
    right sided chemosis | 0
    flexible nasendoscopy made difficult due to thick green secretions | 0
    laboratory tests revealed raised CRP (335 mg/L) | 0
    raised white cell count (24.7 ×10^9/L) | 0
    raised neutrophil count (22.2 ×10^9/L) | 0
    low lymphocyte count (0.5 ×10^9/L) | 0
    raised lactate (2.8 mmol/L) | 0
    pus aspirates collected from both nasal cavities | 0
    microscopy, culture, and sensitivity testing | 0
    Streptococcus pneumoniae isolated | 0
    no evidence of fungal infection | 0
    contrast-enhanced CT of head and sinuses | 1
    CT demonstrated opacification of paranasal sinuses | 1
    bony erosion of lateral walls of both ethmoid sinuses | 1
    soft tissue bulging into right orbit | 1
    bilateral proptosis | 1
    no intracranial abnormality | 1
    patient became increasingly combative | 2
    confused | 2
    aversion to light | 2
    lumbar puncture performed | 3
    pale cloudy fluid macroscopically | 3
    extremely cellular specimen composed mainly of neutrophils | 3
    protein was high (4.07 g/L) | 3
    glucose was low (<0.5 mmol/L) | 3
    Streptococcus pneumoniae isolated | 3
    no evidence of fungal infection | 3
    treatment for sepsis initiated | 4
    treatment for presumed meningitis initiated | 4
    intravenous ceftriaxone | 4
    fluticasone nasal spray | 4
    xylometazoline hydrochloride nasal spray | 4
    regular saline nasal irrigation | 4
    admitted to critical care unit | 4
    joint care of ENT, medical, and critical care teams | 4
    on evening of admission, worsening neurological symptoms | 5
    intubated | 5
    ventilated | 5
    successfully extubated after 8 days | 192
    completed 10-day course of intravenous antibiotics | 240
    discharged home 13 days after admission | 312
    ongoing input from physiotherapy | 312
    occupational therapy teams due to physical deconditioning | 312
    outpatient follow-up with critical care team | 312
    ENT teams arranged | 312
    prescribed 2-week course of betamethasone nasal drops | 312
    6-week course of fluticasone nasal spray | 312
    regular saline nasal irrigation throughout | 312
    3-month follow-up recovering well | 8760
    returned to work full time | 8760
    vivid memories of stay on CCU | 8760
    no signs of post-traumatic stress disorder | 8760
    continued management for CRS with nasal polyposis | 8760
    no further sinus surgery | 8760
    6-month follow-up contrast-enhanced MRI of brain | 4344
    MRI revealed extensive bilateral ethmoid polyposis | 4344
    polyposis extending into maxillary sinuses | 4344
    preseptal space of right orbit | 4344
    hypertrophied inferior turbinates | 4344
    obliterating postnasal space | 4344
    left sided smooth dural enhancement | 4344
    meningeal inflammation | 4344
    Aspergillus specific IgE levels within normal range | 4344
    Alternaria specific IgE levels within normal range | 4344
    <|eot_id|>
    