65 years old | 0
male | 0
admitted to the hospital | 0
abdominal pain | -168
abdominal distension | -168
obstipation | -168
discoloration of abdominal skin | -168
liposuction of the abdomen | -168
gastric bypass | -6048
tachycardia | 0
tachypnoea | 0
normal blood pressure | 0
subcutaneous emphysema of abdominal skin | 0
blackish discoloration of the abdominal skin | 0
erythema | 0
diffuse tenderness | 0
contrast CT scan of the abdomen | 0
hold up of the contrast in the small intestine | 0
dilated jejunum and proximal ileal loops | 0
specks of air in the abdomen | 0
exploratory laparotomy | 24
excision of dead necrotic abdominal skin and subcutaneous tissue | 24
copious amount of seropurulent fluid in the perifascial planes | 24
kinked mid ileal loop | 24
obstruction relieved | 24
perforation in the mid jejunum | 24
perforation repair | 24
debridement | 24
linea alba closed with no. 1 loop nylon | 24
IV fluids | 24
nasogastric aspiration | 24
total parenteral nutrition | 24
altered sensorium | 48
hyponatremia | 48
sepsis | 48
pneumonia | 48
IV antibiotics | 48
E. Coli | 48
Enterococcus | 48
Acticoat dressings | 48
improved wound condition | 336
granulations appeared | 336
reduced soakage | 336
allograft application | 336
reduced exudate | 360
autologous skin grafting | 672
incisional hernia | 8760
incisional hernia repair | 8760