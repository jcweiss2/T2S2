33 years old | 0
female | 0
admitted to the hospital | 0
fever | -210
chills | -210
contact dermatitis | -588
blister on the site of contact dermatitis | -588
antibiotic ointment | -588
steroid ointment | -588
intermittent mild fever | -126
empirical antibiotic treatment | -168
ceftriaxone | -168
azithromycin | -168
discharge | -168
anesthesiology resident | 0
worked in intensive care units | 0
rounded the patients | 0
performed endotracheal intubation | 0
performed central venous catheterization | 0
physical examination | 0
mildly increased white blood cell count | 0
high C-reactive protein | 0
mildly elevated procalcitonin level | 0
normal thyroid function | 0
normal liver function | 0
normal renal function | 0
normal coagulation profile | 0
normal electrolytes | 0
normal lactate levels | 0
polymerase chain reaction results normal | 0
abdominal ultrasonography | 0
obstetric ultrasonography | 0
abdominal and pelvic magnetic resonance imaging scan | 0
S. marcescens cultured in the blood | 48
chorionic tissue infection | 48
empirical cefepime | 0
ceftriaxone | 48
fever again | 96
antibiotic stepped up to cefepime | 96
watery discharge | 552
preterm premature rupture of the membrane | 552
PPROM diagnosed | 552
labor induced | 552
delivered a dead male fetus | 552
IV cefepime | 552
PO clarithromycin | 552
afebrile | 631
leukocytosis normalized | 631
CRP level normalized | 631
discharged | 631
tissue culture from the placenta grew S. marcescens | 631
chorioamnionitis | 631
focal infarct | 631
massive infiltration of neutrophils | 631
spontaneous abortion | 552