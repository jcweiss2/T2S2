80 years old | 0
woman | 0
admitted to the institution via the emergency room | 0
right femur fracture | 0
5-year history of hypertension | -43800
hypertension | -43800
medication regimen of an antihypertensive agent | -43800
aspirin | -43800
obesity | 0
depression | 0
delirium symptoms | 0
brain CT | 0
severe stenosis of the middle cerebral artery (MCA) | 0
old localized infarction of the basal ganglia | 0
diffuse atrophy of the brain | 0
cardiomegaly | 0
1 degree A-V block | 0
ejection fraction of 65% | 0
preoperative PT/PTT was 12.7/24.4 seconds | 0
INR was 1.15 | 0
pH 7.376 | 0
PaO2 78.6 mmHg | 0
PaCO2 27.5 mmHg | 0
total hip replacement surgery scheduled | 96
aspirin maintained until the 3rd hospital day | 72
standard monitoring devices applied | 96
left radial artery cannulated | 96
BP 140/70 mmHg | 96
heart rate 80 beats/min | 96
O2 saturation 98% | 96
spinal anesthesia administered | 96
right lateral position | 96
L3-4 interspace | 96
0.5% hyperbaric bupivacaine 8 mg | 96
supine position | 96
unresponsive | 96
BP 70/40 mmHg | 96
HR 40-45 beats/min | 96
ephedrine administration | 96
epinephrine 10 µg | 96
crystalloid infusion | 96
endotracheal intubation | 96
manual ventilation | 96
norepinephrine 0.1 µg/kg/min | 96
dopamine 2 µg/kg/min | 96
BP 60/40 mmHg | 96
HR 110 beats/min | 96
IV epinephrine 0.02 µg/kg/min | 96
PaO2 488.9 mmHg | 96
PaCO2 30.8 mmHg | 96
FiO2 1.0 | 96
EtCO2 28 mmHg | 96
O2 saturation 99% | 96
high spinal anesthesia suspected | 96
central venous catheterization | 96
right internal jugular vein | 96
central venous pressure 30 mmHg | 96
TEE performed | 96
right atrium (RA) enlargement | 96
right ventricle (RV) enlargement | 96
straightening of the interventricular septum | 96
hypokinesia | 96
PE diagnosis | 96
IV heparin 5,000 IU | 96
heparin maintained at 1,000 IU/hr | 96
milrinone 50 µg/kg | 96
milrinone maintained at 0.5 µg/kg/min | 96
pH 7.224 | 96
PaO2 55.2 mmHg | 96
PaCO2 52.8 mmHg | 96
operation postponed | 96
transported to ICU | 96
heart rate decreased to 30 beats/min | 96
cardiopulmonary resuscitation | 96
chest 3D PTCA | 96
non-contrast brain CT | 96
low density ovoid thromboembolism | 96
enlargement of right atrium and ventricle | 96
low density large acute infarct | 96
gyral swelling of the right insula and temporal lobe | 96
heart rate decreased to 30 beats/min | 113
resuscitation ineffective | 113
died | 113
PaCO2 27.5 mmHg |7 0
