68 years old | 0
    male | 0
    type II diabetes mellitus | 0
    peripheral neuropathy | 0
    hypertension | 0
    chronic obstructive pulmonary disease | 0
    home oxygen | 0
    bipolar depression | 0
    gastroesophageal reflux | 0
    shortness of breath | -336
    cough | -336
    decrease in exercise tolerance | -336
    intermittent diarrhea | -336
    treated with vancomycin | 0
    treated with piperacillin/tazobactam | 0
    transferred to medical intensive care unit | 0
    dopamine started | 0
    hypotension | 0
    presumed sepsis | 0
    condition stabilized | 0
    transferred to medical floor | 0
    pulmonary embolus | 0
    colonic distension | 0
    profuse watery diarrhea | 0
    colonic pseudo-obstruction (Ogilvie's syndrome) | 0
    nasogastric tube placed | 0
    rectal tube placed | 0
    renal service consulted | 0
    hypokalemia | 0
    difficult to control with potassium supplementation | 0
    aspirin 81 mg daily | 0
    atorvastatin 80 mg daily | 0
    budesonide/formoterol | 0
    levalbuterol | 0
    tiotroprium | 0
    insulin | 0
    pantoprazole 40 mg daily |?0
    piperacillin/tazobactam | 0
    potassium chloride 100 mEq daily | 0
    blood pressure 103/50 mm Hg | 0
    pulse 102 beats per minute | 0
    respiratory rate 24 breaths per minute | 0
    tachypneic | 0
    using accessory muscles | 0
    rhonchi in anterior lung fields | 0
    abdomen distended | 0
    hypoactive bowel sounds | 0
    tenderness in right upper quadrant | 0
    tenderness in midepigastric area | 0
    trace lower extremity edema | 0
    Foley catheter in place | 0
    rectal tube in place | 0
    serum sodium 146 mmol/l | 0
    serum chloride 118 mmol/l | 0
    serum potassium 2.7 mmol/l | 0
    serum bicarbonate 19.9 mmol/l | 0
    blood urea nitrogen 6.1 mmol/l | 0
    serum creatinine 110 μmol/l | 0
    serum potassium on admission 4.1 mmol/l | 0
    arterial pH 7.27 | 0
    arterial pCO2 36.9 mm Hg | 0
    arterial bicarbonate 17.1 mEq/l | 0
    urine sodium 49 mmol/l | 0
    urine potassium 20 mmol/l | 0
    urine chloride 90 mmol/l | 0
    urine anion gap -21 | 0
    24-hour urine potassium 9.1 mmol | 0
    stool sodium <10 mmol/l | 0
    stool potassium 139.7 mmol/l | 0
    colonic distension (13 cm) | 0
    diagnosis of severe gastrointestinal potassium wasting | 0
    received potassium chloride >100 mmol/day | 0
    serum potassium 3.5–4.0 mmol/l | 0
    respiratory status deteriorated | 0
    family withdrew care | 0
    patient expired | 0

    68 years old | 0
    male | 0
    type II diabetes mellitus | 0
    peripheral neuropathy | 0
    hypertension | 0
    chronic obstructive pulmonary disease | 0
    home oxygen | 0
    bipolar depression | 0
    gastroesophageal reflux | 0
    shortness of breath | -336
    cough | -336
    decrease in exercise tolerance | -336
    intermittent diarrhea | -336
    treated with vancomycin | 0
    treated with piperacillin/tazobactam | 0
    transferred to medical intensive care unit | 0
    dopamine started | 0
    hypotension | 0
    presumed sepsis | 0
    condition stabilized | 0
    transferred to medical floor | 0
    pulmonary embolus | 0
    colonic distension | 0
    profuse watery diarrhea | 0
    colonic pseudo-obstruction (Ogilvie's syndrome) | 0
    nasogastric tube placed | 0
    rectal tube placed | 0
    renal service consulted | 0
    hypokalemia | 0
    difficult to control with potassium supplementation | 0
    aspirin 81 mg daily | 0
    atorvastatin 80 mg daily | 0
    budesonide/formoterol | 0
    levalbuterol | 0
    tiotroprium | 0
    insulin | 0
    pantoprazole 40 mg daily | 0
    piperacillin/tazobactam | 0
    potassium chloride 100 mEq daily | 0
    blood pressure 103/50 mm Hg | 0
    pulse 102 beats per minute | 0
    respiratory rate 24 breaths per minute | 0
    tachypneic | 0
    using accessory muscles | 0
    rhonchi in anterior lung fields | 0
    abdomen distended | 0
    hypoactive bowel sounds | 0
    tenderness in right upper quadrant | 0
    tenderness in midepigastric area | 0
    trace lower extremity edema | 0
    Foley catheter in place | 0
    rectal tube in place | 0
    serum sodium 146 mmol/l | 0
    serum chloride 118 mmol/l | 0
    serum potassium 2.7 mmol/l | 0
    serum bicarbonate 19.9 mmol/l | 0
    blood urea nitrogen 6.1 mmol/l | 0
    serum creatinine 110 μmol/l | 0
    serum potassium on admission 4.1 mmol/l | 0
    arterial pH 7.27 | 0
    arterial pCO2 36.9 mm Hg | 0
    arterial bicarbonate 17.1 mEq/l | 0
    urine sodium 49 mmol/l | 0
    urine potassium 20 mmol/l | 0
    urine chloride 90 mmol/l | 0
    urine anion gap -21 | 0
    24-hour urine potassium 9.1 mmol | 0
    stool sodium <10 mmol/l | 0
    stool potassium 139.7 mmol/l | 0
    colonic distension (13 cm) | 0
    diagnosis of severe gastrointestinal potassium wasting | 0
    received potassium chloride >100 mmol/day | 0
    serum potassium 3.5–4.0 mmol/l | 0
    respiratory status deteriorated | 0
    family withdrew care | 0
    patient expired | 0