88 years old | 0
hypertension | -720
atrial fibrillation | -720
unstable angina | -720
left-side motor weakness | 0
right-side eyeball deviation | 0
admitted to a district hospital | 0
right middle cerebral artery infarction | 0
tissue plasminogen activator | 0
dyspnea | 168
unstable vital signs | 168
blood pressure 80/40 mmHg | 168
heart rate 150 beats/min | 168
respiration 44 breaths/min | 168
body temperature 39.1℃ | 168
O2 saturation 94% | 168
septic shock | 168
intubated | 168
left subclavian venous catheterization attempted | 168
lidocaine injected | 168
left subclavian vein identified | 168
Seldinger-type central venous catheter set used | 168
guidewire passed through introducer needle | 168
minimal resistance encountered during guidewire insertion | 168
guidewire advanced approximately 30 cm | 168
guidewire could not be advanced further | 168
attempts to withdraw guidewire failed | 168
chest X-ray showed guidewire knotted and kinked | 168
transferred to our hospital | 168
portable chest X-ray performed | 0
subclavian venogram performed | 0
X-ray revealed guidewire knotted and kinked | 0
guidewire folded back and entered mediastinum | 0
subclavian venogram revealed guidewire not perforated subclavian vein | 0
guidewire knotted, kinked, and extended extravascularly | 0
subclavian vein intact | 0
surgical exploration decided | 0
general anesthesia | 0
initial vital signs: blood pressure 100/50 mmHg | 0
initial heart rate 134 beats/min | 0
initial respiration 25 breaths/min | 0
initial O2 saturation 96% | 0
anesthesia induced with etomidate | 0
anesthesia induced with rocuronium | 0
noninvasive blood pressure cuff applied on right arm | 0
arterial catheter placed in left radial artery | 0
femoral venous catheter applied at left femoral vein | 0
7-cm incision made | 0
guidewire beneath subclavian vein | 0
tangled part of wire kinked between sternocleidomastoid muscles | 0
vessels not damaged | 0
guidewire cut to untangle | 0
guidewire pulled out from mediastinum | 0
entire guidewire removed | 0
postoperative intensive care unit | 24
discharged to ward | 48
