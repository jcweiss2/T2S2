61 years old | 0
male | 0
admitted to hospital | 0
sepsis | 0
Candida albicans | 0
hypertension | -672
dyslipidemia | -672
type 2 diabetes | -672
urinary retention | -672
phimosis | -672
balanitis xerotica obliterans | -672
urethral strictures | -672
aspirin | -672
bisoprolol | -672
ezetimibe | -672
empagliflozin | -672
gliclazide | -672
metformin | -672
ramipril | -672
vomiting | -336
fever | -336
flank pain | -336
pyelonephritis | -336
left hydronephrosis | -336
left nephrostomy tube | -336
hypoxia | -336
pulmonary edema | -336
fluconazole | -336
caspofungin | -336
vision loss | 0
Code Stroke | 0
CT/CTA | 0
hemoglobin 103 g/L | 0
C-reactive protein 47.3 mg/L | 0
sedimentation rate 75 mm/h | 0
visual acuity 20/20 OD | 0
visual acuity NLP OS | 0
RAPD | 0
mild right optic disc edema | 0
cotton wool spots | 0
left pallid optic disc edema | 0
OCT | 0
increased thickness 127 μm OD | 0
blood pressure 98/40 | -1
diagnosis of anterior ischemic optic neuropathy | 0
blood pressure medications held | 0
salt tablets | 0
midodrine | 0
hydration | 0
blood pressure improved | 24
visual function stabilized | 24
optic disc edema improved | 720
OCT retinal nerve fiber layer resolved | 720
visual acuity 20/20 OD | 720
visual acuity NLP OS | 720
Humphrey visual fields | 720
sepsis-induced NAION | 0
hypotension | -1
anemia | 0
disk-at-risk appearance | -672
vascular risk factors | -672
bilateral optic disc edema | 0
increased intracranial pressure | 0
hypertensive crisis | 0
infection/inflammation | 0
toxic/nutritional conditions | 0
demyelinating conditions | 0
broad differential diagnosis | 0
early recognition | 0
aggressive blood pressure control | 0
partial visual recovery | 720