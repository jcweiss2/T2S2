63 years old | 0
male | 0
achalasia | 0
dyspepsia | 0
referred to the hospital | 0
sudden onset | 0
severe right chest pain | 0
epigastric pain | 0
chest retrosternal pain |'0
respiratory distress | 0
tachycardic | 0
arterial pressure | 0
no fever | 0
diminished breath sounds | 0
pain | 0
tenderness of epigastric | 0
normal laboratory findings | 0
O2 saturation | 0
computed tomography scan | 0
pneumomediastinum | 0
pleural effusion | 0
collapsed right lobe of the lung | 0
Candida albicans in pleural space | 0
extravasation to the right pleural space | 0
esophageal content in pleural space | 0
general condition worsened | 0
admitted to ICU | 0
intubated | 0
antibiotics | 0
chest physical therapy | 0
intravenous fluids | 0
nasogastric tube feeding | 0
WBC count elevated | 72
BUN elevated | 72
potassium elevated | 72
tachyarrhythmia | 72
multiple organ failures | 96
kidney failure | 96
hemodialysis | 96
kidney function normalized | 96
thoracotomy | 96
continuation of sepsis | 96
accumulation of pus | 96
secretion of the right pleural space | 96
longitudinal rupture in upper esophagus | 96
patient unstable | 96
noradrenaline | 96
vasopressin | 96
T-tube implanted | 96
sutures | 96
chest tubes inserted | 96
ventilator support | 96
vasopressor | 96
piperacillin/tazobactam | 96
esophageal stents placed | 96
oral liquid feeding | 120
ICU stay | 936
discharged from hospital | 1008
tracheostomy | 240
follow-up after two months | 1824
