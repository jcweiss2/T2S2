45 years old | 0
female | 0
admitted to the hospital | 0
pain in abdomen | -48
vomiting | -48
caesarean section delivery | -52560
incisional hernia | -4032
laparoscopic incisional hernia repair | -4032
ePTFE mesh placed intraperitoneally | -4032
tackers | -4032
trans-abdominal polypropylene sutures | -4032
vomiting on and off | -2688
conscious | 0
oriented | 0
pulse rate 120/min | 0
blood pressure 50 mmHg systolic | 0
added sounds on chest auscultation | 0
mild distension | 0
tenderness | 0
rigidity | 0
guarding | 0
7cm fluctuant swelling in right lumbar quadrant | 0
blackish discoloration of overlying skin | 0
Hb 7.5 g/dl | 0
Total Leucocyte Count 5840 cells/cmm | 0
blood glucose 66 mg/dl | 0
serum creatinine 1.4 mg/dl | 0
serum albumin 1.3 g/dl | 0
serum sodium 142.6 meq/l | 0
serum potassium 3.1 meq/l | 0
ultrasonography abdomen loculated collection in pelvis (~60cc) | 0
parietal wall collection (~100cc) in right lower abdomen | 0
communicating with peritoneal cavity | 0
scar dehiscence | 0
X-ray chest patchy-confluent consolidation in bilateral lung fields | 0
admitted to ICU | 0
intravenous fluids | 0
inotropic drugs | 0
ventilatory support | 0
difficulty in respiration | 0
falling arterial oxygen saturation | 0
operated | 0
necrotising fasciitis of overlying abdominal wall | 0
infected mesh densely adhered to gut | 0
feculent fluid | 0
dense cohesive adhesions | 0
two nearby small bowel perforations | 0
liberal debridement of overlying anterior abdominal wall | 0
maximum resection of implanted mesh | 0
small bowel segmental resection | 0
exteriorisation of bowel ends | 0
multiorgan dysfunction syndrome | 72
expired | 72
