45 years old | 0
male | 0
admitted to the emergency department | 0
fever | -144
temperature 39°C | -144
cough | -144
dyspnoea | -144
diarrhoea | -144
vomiting | -144
abdominal pain | -144
bilateral crackles on lung bases | 0
severe pain in epigastrium | 0
rigidity of abdominal wall | 0
guarding of abdominal wall | 0
SpO2 82% | 0
heart rate 109 beats per minute | 0
blood pressure 89/47 mmHg |%0
intubated | 0
mechanically ventilated | 0
resuscitated | 0
low-dose noradrenaline | 0
crystalloid fluids | 0
SARS-CoV-2 positive | 0
leukocytosis 20×10³ white blood cells | 0
lymphocytopenia 0.47×10³/L | 0
increased C-reactive protein 99 mg/L | 0
increased lactate dehydrogenase 997 U/L | 0
increased lactate 6 mmol/L | 0
increased d-dimers 4.1 μg/mL | 0
blood urea nitrogen 6.1 mmol/L | 0
creatinine 119 μmol/L | 0
chest CT bilateral peripheral ground-glass opacities | 0
infiltrates | 0
pulmonary embolism | 0
abdominal CT thickened bowel wall | 0
portal vein thrombosis | 0
duplex ultrasonography excluded deep vein thrombosis | 0
emergency exploratory laparotomy | 24
contained small intestinal perforation | 24
peritonitis | 24
resection of ischaemic jejunum | 24
epithelial necrosis | 24
haemorrhagic infarction | 24
neutrophilic inflammation | 24
fibrin deposition within lamina propria | 24
admitted to ICU | 24
ribavirin 400 mg every 12 hours | 24
meropenem 0.5 g intravenously every 12 hours | 24
vancomycin 15 mg/kg loading dose | 24
therapeutic anticoagulation enoxaparin 75 mg | 24
ARDS-net ventilation | 24
hydrocortisone | 24
vasopressors | 24
supportive ICU care | 24
acute kidney injury (AKI) | 24
blood urea nitrogen 7.9 mmol/L | 24
creatinine 309 μmol/L | 24
mild metabolic acidosis | 24
hyperkalaemia | 24
anuric | 24
shock necessitating vasopressors | 24
continuous renal replacement therapy (CRRT) | 24
CytoSorb filter | 24
transfusion two packs red blood cells | 24
diuresis initiated | 72
weaned off vasopressors | 72
lactate normalized | 72
inflammatory biomarkers normalized | 72
CRRT discontinued | 72
oxygenation improved | 72
PaO2/FiO2 ratio >300 | 168
extubated | 168
renal function normalized | 336
broad-spectrum antibiotics | 336
therapeutic anticoagulation continued | 336
RT-PCR negative for COVID-19 | 456
lupus anticoagulant negative | 576
antiphospholipid antibodies negative | 576
antineutrophil cytoplasmic antibodies negative | 576
thrombophilia screening negative | 576
blood cultures negative | 576
urine cultures negative | 576
sputum cultures negative | 576
discharged | 816
oral rivaroxaban prescribed | 816
