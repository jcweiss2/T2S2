19 years old | 0
female | 0
admitted to the hospital | 0
vaginal bleeding | -216
fresh blood and clots | -216
vaginal bleeding started | -216
vaginal bleeding persisted | -9
vesicle-like tissue present | -24
married | -8760
spontaneous full-term singleton birth | -7300
antenatal visit | -168
referred to obstetrician | -168
ultrasound screening | -168
suspicious for molar pregnancy | -168
referred to hospital | -168
curettage planned | 0
vital signs normal | 0
physical examination | 0
speculum examination | 0
insignificant bleeding | 0
no mass infiltration | 0
anemia | 0
leukocytes 9630/uL | 0
platelets 396 000/µL | 0
β-hCG level 1000×103 mIU/mL | 0
thyroid function normal | 0
chest X-rays normal | 0
ultrasound scan | 0
enlarged uterus | 0
vesicular appearance | 0
suspected molar pregnancy | 0
blood transfusion | 0
vacuum curettage | 120
mass on left labia minora | 120
mass measured 3×3×2 cm | 120
suspected hematoma | 120
additional sharp curettage | 120
uterine cavity completely removed | 120
conservative management | 120
pain in genital area | 124
vital signs deteriorated | 124
went into shock | 124
vulvar mass | 124
perforation | 124
active bleeding | 124
emergency evacuation | 124
hematoma incised | 124
blood and clot evacuated | 124
vesicle-like tissue found | 124
fragile tissue found | 124
bleeding controlled | 124
suspected stage II GTN | 124
histopathological examination | 124
chronic villi with cystic dilatation | 124
hydrophilic avascular degeneration | 124
cytotrophoblasts and syncytiotrophoblasts | 124
excessive proliferation | 124
nuclei within normal limits | 124
blood clot in decidua | 124
no malignant tumor cells | 124
final histopathologic diagnosis | 124
complete mole with excessive trophoblastic cell proliferation | 124
reevaluation of histopathologic examination | 124
partial hydatidiform mole | 124
immunohistochemical examination | 124
p53 positive | 124
transferred to ICU | 124
oxygen saturation 80% | 124
prolonged intubation | 124
hypoxia | 124
postoperative hemoglobin 2.3 g/dL | 124
transfusion | 124
hemoglobin 9 g/dL | 124
bilateral pneumonia | 148
leukocytosis | 148
sepsis | 148
antibiotics | 148
pulmonary edema | 196
metabolic encephalopathy | 196
died due to sepsis | 528
cause of death unknown | 528
refused autopsy | 528