55 years old | 0
male | 0
road traffic accident | -2
multiple tissue injuries | -2
loss of consciousness | -2
right lobe liver injury | -2
subarachnoid hemorrhages | -2
multiple contusions | -2
admitted to emergency department | 0
high-grade fever | 48
sepsis | 48
total leukocyte count increased | 48
erythrocyte sedimentation rate increased | 48
blood culture showed growth of smooth, nonpigmented mucoid colonies | 48
Gram-positive cocci in clusters | 48
catalase positive | 48
negative for tube coagulase | 48
negative for mannitol fermentation | 48
negative for ornithine decarboxylase | 48
identified as S. haemolyticus | 48
resistance to penicillin | 48
resistance to cefoxitin | 48
resistance to gentamicin | 48
resistance to erythromycin | 48
resistance to clindamycin | 48
vancomycin sensitive | 48
LZ resistant | 48
cfr gene detected | 48
treated with vancomycin | 72
died of infection | 120
mucoid variant of S. haemolyticus | 48
capsular polysaccharides production | 48
enhanced virulence | 48
LZ resistance without exposure to LZ | 48
mucoid colonies indistinguishable from Klebsiella spp. | 48
retained mucoid characteristic on serial subcultures | 72
higher virulence of the mucoid strain | 120
comorbidities in the patient | 120