history of difficult-to-manage bronchial asthma | -720
hospitalized for acute exacerbations | -720
dry cough | -24
progressive dyspnea | -24
psychomotor agitation | -24
audible wheezing | -24
admitted in critical condition | 0
diaphoretic | 0
tachycardic | 0
dyspneic | 0
supraclavicular retractions | 0
respiratory rate of 30 breaths/minute | 0
ambient oxygen saturation 87% | 0
auscultation with abolished vesicular murmur | 0
Glasgow coma scale 12/15 | 0
arterial blood gases analysis | 0
respiratory acidosis | 0
hypoxemia | 0
invasive ventilatory support | 0
midazolam administration | 0
propofol administration | 0
hydrocortisone administration | 0
magnesium sulfate administration | 0
antibiotics administration | 0
neuromuscular blocking agents administration | 48
improvement in ABG | 96
ventilatory weaning | 96
suspension of dual sedation | 96
suspension of NMB | 96
light sedation with dexmedetomidine | 96
weakness of the neck flexor muscles | 144
facial paresis | 144
quadriplegia | 144
flaccid hyporeflexia | 144
preserved sensitivity | 144
normal cranial nerves | 144
brain and cervical MRI | 144
cerebrospinal fluid study | 144
MRC score 37 points | 144
electromyography | 144
denervation and irritability | 144
polyneuropathic compromise | 144
axonal pattern in conduction velocity | 144
diagnosis of ICUAW | 144
physiotherapy | 144
comprehensive rehabilitation | 144
ventilator withdrawal | 240
hospital discharge | 720
MRC score 55 points | 720
normal ABG control | 720
symptomatic resolution | 720