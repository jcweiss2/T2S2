38 years old|0
male|0
presented to the emergency department|0
fever|0
cough|0
shortness of breath|0
myalgia|0
BMI of 29.9|0
history of daily vaping|0
no history of recent travel|0
no known contact with COVID-19 positive individuals|0
CT angiogram|0
no pulmonary embolism|0
bilateral numerous multifocal ground glass opacities|0
multifocal viral pneumonia|0
SARS COV2 PCR nasopharyngeal swab test|0
confirmed COVID-19 positive|0
placed on droplet precautions|0
contact isolation|0
blood culture|0
sputum culture|0
urine legionella testing|0
sputum legionella testing|0
mycoplasma IGM tests|0
negative results|0
subcutaneous Heparin|0
D-dimer elevated|0
decompensated|120
intubated|120
acute hypoxemic respiratory failure|120
admitted to the intensive care unit|120
placed on Plaquenil|120
supplemental oxygen|120
albuterol sulfate|120
tiotropium bromide|120
Tocilizumab|120
Zithromax|120
acute renal failure|144
sepsis|816
toxic metabolic encephalopathy|936
temperature 100°F|0
pulse 122|0
blood pressure 141/81|0
white blood cell low|0
red blood cell normal|0
platelet high|0
neutrophil percentage high|0
lymphocyte percentage high|0
C-reactive protein high|0
creatinine high|0
PTT high|0
fibrinogen high|0
pro-calcitonin high|0
lactate dehydrogenase high|0
alanine aminotransferase high|0
aspartate aminotransferase high|0
calcium low|24
potassium high|24
glucose high|24
insulin therapy|24
continuous veno-venous hemofiltration|24
intermittent hemodialysis|24
troponin-I high|240
creatinine kinase high|240
creatinine kinase maximum|408
anemia|1104
hemoglobin 6.8|1104
transfused|1104
Hemophagocytic lymphohistiocytosis syndrome|1104
delirium|1104
toxic metabolic encephalopathy|1104
prolonged hospitalization|1104
infections|1104
CT chest scan|1104
persistent bilateral posterior thoracic and shoulder muscular findings|1104
magnetic resonance cholangiopancreatography|1464
elevated alkaline phosphatase|1464
no abnormalities in pelvic and proximal thigh muscles|1464
interdisciplinary rehabilitation therapy program|2160
discharge arrangements being made|2160
