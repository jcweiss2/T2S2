57 years old | 0
male | 0
smoking history | 0
admitted to the hospital | 0
fever | -48
cough | -48
sputum | -48
dyspnea | -24
hypothermia | 0
tachypnea | 0
hypoxemia | 0
tachycardia | 0
low blood pressure | 0
moist rale | 0
hypoxygen | 0
metabolic acidosis | 0
hyperlactatemia | 0
infection | 0
multiple organ injury | 0
lung consolidation | 0
fluid resuscitation | 0
continuous renal replacement treatment | 0
organ protective therapy | 0
empiric antibiotic therapy | 0
piperacillin tazobactam | 0
moxifloxacin | 0
nasal intubation | 0
mechanical ventilation | 0
prone position ventilation | 0
Klebsiella pneumoniae | 72
antimicrobial susceptibility testing | 72
hvKP | 72
string test | 72
wax moth larvae test | 72
hypoxemia improved | 72
unstable hemodynamics | 72
norepinephrine | 72
thoracic CT | 240
lung abscess | 240
CEUS | 288
contrast-enhanced ultrasound | 288
SonoVue | 288
CEUS-guided drainage | 288
pigtail tube | 288
hypoxemia improved | 384
hemodynamics improved | 384
weaned from ventilator | 384
thoracic CT | 504
lung lesion improved | 504