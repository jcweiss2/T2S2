74 years old | 0
female | 0
Hispanic | 0
from Ecuador | 0
type 2 diabetes mellitus | -672
fever | -120
jaundice | -120
right upper quadrant abdominal pain | -120
unintentional weight loss | -720
vomiting | -120
denies chest pain | -120
denies dyspnea | -120
denies melena | -120
denies hematochezia | -120
denies dysuria | -120
denies hematuria | -120
no history of cigarette | 0
no history of alcohol | 0
no history of substance abuse | 0
no family history of cancer | 0
elevated serum alkaline phosphatase | 0
serum creatinine of 3.83 mg/dL | 0
international normalized ratio (INR) of 1.4 | 0
serum lactate dehydrogenase (LDH) of 471 U/L | 0
leukocytosis | 0
monocytosis | 0
thrombocytopenia | 0
macrocytic anemia | 0
hemoglobin (Hb) 9 g/dL | 0
mean corpuscular volume (MCV) of 102.4 fL | 0
no blasts identified | 0
admitted to the ICU | 0
treated with broad-spectrum antibiotics | 0
cholelithiasis | 0
thickened gallbladder wall | 0
positive sonographic Murphy sign | 0
dilated common bile duct | 0
endoscopic retrograde cholangiopancreatography (ERCP) | 24
purulence in the common bile duct | 24
stone in the common bile duct | 24
stone removed | 24
plastic stent placed in the common bile duct | 24
laparoscopic cholecystectomy | 48
insertion of a Jackson-Pratt drain | 48
gangrenous gallbladder | 48
given crystalloid fluid | 48
given platelets | 48
given irradiated packed red blood cells (PRBCs) | 48
continued fever | 72
progressive leukocytosis | 72
sepsis | 72
active treatment discontinued | 96
made as comfortable as possible | 96
histopathology of the gallbladder | 120
myeloblasts in the gallbladder | 120
promyelocytes in the gallbladder | 120
myelocytes in the gallbladder | 120
immunohistochemistry | 120
neoplastic cells positive for lysozyme | 120
neoplastic cells positive for CD68 | 120
neoplastic cells positive for CD33 | 120
neoplastic cells positive for HLA-DR | 120
neoplastic cells positive for CD117 | 120
neoplastic cells positive for myeloperoxidase | 120
neoplastic cells positive for CD56 | 120
neoplastic cells negative for CD34 | 120
granulocytic sarcoma | 120
extramedullary acute myelomonocytic leukemia (AML M5) | 120
death | 168