33 years old | 0
female | 0
admitted to the emergency department | 0
cardiac arrest | 0
liposuction of thighs | -0.75
harvesting 1.5 L of fat | -0.75
somnolent | -0.25
stable vital signs | -0.25
blood pressure 170/90 mmHg | -0.25
suspected hypoglycemia | -0.25
administered oral dextrose solution | -0.25
no improvement | -0.25
dizzy | 2
rapid decline of mental status | 2
tonic-clonic seizure | 2
loss of consciousness | 2
gasping | 2.25
cyanotic | 2.25
drooling | 2.25
cardiopulmonary arrest | 2.25
resuscitation | 2.25
asystole | 2.5
intubated | 2.5
resuscitation | 2.5
return of spontaneous circulation | 2.5
power-assisted liposuction technique | -0.75
use of five vials of 50 mL lidocaine 2% | -0.75
total dose of lidocaine 5000 mg | -0.75
prior use of same procedure and anesthesia | -2160
abdominal liposuction | -2160
normal sinus rhythm | 2.5
no QT prolongation | 2.5
QTc 466 ms | 2.5
normal QRS interval 100 ms | 2.5
no ST- or T-wave abnormalities | 2.5
Glasgow Coma Scale 3T | 2.5
pupils equal in size bilaterally | 2.5
reactive to light | 2.5
preserved corneal and oculocephalic reflexes | 2.5
downward Babinski reflex bilaterally | 2.5
arterial blood gas analysis | 2.5
pH 7.34 | 2.5
CO2 pressure 39.9 mmHg | 2.5
O2 pressure 131 mmHg | 2.5
bicarbonate concentration 20.8 mmol/L | 2.5
white blood cell count 9.8 × 10^9/L | 2.5
polymorphonuclear cells 41% | 2.5
hemoglobin level 10.4 g/dL | 2.5
platelet count 336 × 10^6/L | 2.5
troponin 0.003 ng/mL | 2.5
sodium concentration 144 mmol/L | 2.5
potassium 3.5 mmol/L | 2.5
chloride 99 mmol/L | 2.5
bicarbonate 16 mmol/L | 2.5
glucose 346 mg/dL | 2.5
blood urea nitrogen 13 mg/dL | 2.5
creatinine 1.0 mg/dL | 2.5
aspartate aminotransferase 225 IU/L | 2.5
alanine aminotransferase 238 IU/L | 2.5
γ-glutamyl transpeptidase 12 IU/L | 2.5
alkaline phosphatase 55 IU/L | 2.5
lactate 17.55 mmol/L | 2.5
serum lidocaine level 5.30 µg/mL | 2.5
CT scan of brain | 2.5
CT angiography of chest | 2.5
bilateral consolidations | 2.5
aspiration pneumonitis | 2.5
no intracranial bleeding | 2.5
no pulmonary embolism | 2.5
no aortic dissection | 2.5
antibiotic therapy | 2.5
generalized myoclonic jerks | 2.5
anoxic brain injury | 2.5
valproic acid | 2.5
admitted to intensive care unit | 2.5
magnetic resonance imaging of brain | 72
severe hypoxic-ischemic brain injury | 72
electroencephalogram | 72
electrocerebral silence | 72
increase in brain edema and pressure | 120
electrolytes disturbances | 120
multiple nosocomial infections | 120
end-organ damage | 120
septic shock | 1440
death | 1440