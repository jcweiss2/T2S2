67 years old | 0  
    male | 0  
    severe rheumatoid arthritis | 0  
    tocilizumab | 0  
    dyspnea | 0  
    chest pain | 0  
    tachycardia | 0  
    tachypnea | 0  
    hypotension | 0  
    elevated WBC count (48.6 × 103/uL) | 0  
    lactic acid elevated (8.9 mmol/L) | 0  
    SGOT (AST) elevated (2552) | 0  
    SGPT (ALT) elevated (5198) | 0  
    sinus tachycardia | 0  
    low voltage on electrocardiography | 0  
    emergent intubation | 0  
    pericardiocentesis | 0  
    removal of 800 mL cloudy, milky fluid | 0  
    admitted to ICU | 0  
    provisional diagnosis of rheumatoid pericardial effusion | 0  
    cardiac tamponade | 0  
    septic shock | 0  
    pressor support | 0  
    broad-spectrum antibiotics | 0  
    blood culture negative | 0  
    urine culture negative | 0  
    indium scan showing WBC accumulation in upper abdomen | 0  
    discharge to skilled nursing facility | 0  
    recurrent shortness of breath | 336  
    moderate pericardial effusion | 336  
    pericardial window placement | 336  
    generalized abdominal pain | 336  
    back pain | 336  
    recurrent leukocytosis | 336  
    pericardial fluid lipase elevated (24000 U/L) | 336  
    CT showing gas-containing fluid collection anterior to heart | 336  
    fluid collections in pancreatic head and neck | 336  
    surgical exploration revealing pancreaticopericardial fistula | 336  
    infected pericardial window | 336  
    irrigation of pericardial space | 336  
    drain placement | 336  
    jaundice | 336  
    wound infection | 336  
    enzymatic breakdown of wound | 336  
    wound vacuum placement | 336  
    somatostatin | 336  
    EGD | 336  
    ERCP revealing organized necrosis | 336  
    communication to lumen | 336  
    side branch disruption at head | 336  
    filling of lesser sac | 336  
    stent placement into pancreatic duct | 336  
    hypotension | 336  
    unable to maintain perfusion | 336  
    emergent family meeting | 336  
    decision to limit treatment to comfort measures | 336  
    patient expired | 336  
    acute pancreatitis | 0  
    gallstone-induced pancreatitis excluded | 0  
    ethanol-induced pancreatitis excluded | 0  
    hypertriglyceridemia-induced pancreatitis excluded | 0  
    tocilizumab possible role | 0  
    pancreatic pseudocyst | 0  
    pancreatic necrosis | 0  
    superimposed infection | 336  
    pancreaticopericardial fistula | 336  
    infected pericardial window | 336  

    67 years old | 0  
    male | 0  
    severe rheumatoid arthritis | 0  
    tocilizumab | 0  
    dyspnea | 0  
    chest pain | 0  
    tachycardia | 0  
    tachypnea |D