22 years old | 0
male | 0
admitted to the hospital | 0
mild COVID-19 illness | -72
sore throat | -72
loss of sense of smell | -72
positive COVID-19 PCR | -72
full recovery | -40
resolution of symptoms | -40
negative PCR | -40
first dose of inactivated SARS-CoV-2 vaccine | -30
asymptomatic | -30
second dose of inactivated SARS-CoV-2 vaccine | 0
headache | 2
fatigue | 2
fever | 24
sore throat | 24
abdominal pain | 24
high-grade fever | 96
myalgia | 96
nausea | 96
vomiting | 96
diarrhea | 96
faint erythematous non-itchy rash | 96
dry irritant cough | 96
no shortness of breath | 96
no chest discomfort | 96
no urinary symptoms | 96
no pain or swelling of joints | 96
temperature of 39°C | 96
systolic blood pressure of 110 mm Hg | 96
tachycardia | 96
dry mucous membranes | 96
congested throat | 96
bilateral conjunctival injection | 96
left conjunctival hemorrhage | 96
generalised erythematous maculopapular rash | 96
no enlarged peripheral lymph nodes | 96
no audible cardiac murmurs | 96
clear chest | 96
unremarkable abdomen examination | 96
SARS-CoV-2 PCR negative | 96
SARS-CoV-2 IgG positive | 96
throat swab negative for group A streptococcus | 96
sputum culture showed mixed flora | 96
bacterial blood cultures negative | 96
significant proteinuria | 96
ANA negative | 96
dsDNA negative | 96
c-ANCA negative | 96
p-ANCA negative | 96
C3 reduced | 96
C4 reduced | 96
admitted to ICU | 96
treated with ceftriaxone | 96
treated with levofloxacin | 96
intravenous hydrocortisone | 96
haemodynamic stability | 120
discontinued hydrocortisone | 120
persistent fever | 120
facial puffiness | 120
generalised body oedema | 120
tachycardia | 120
diarrhea | 120
myalgia | 120
anasarca | 120
renal impairment | 120
significant proteinuria | 120
ECG showed sinus tachycardia | 120
non-specific T-wave abnormalities | 120
troponin-I raised | 120
pro-BNP raised | 120
severe tricuspid regurgitation | 120
pulmonary hypertension | 120
moderately dilated right atrium and ventricle | 120
normal systolic function | 120
mildly reduced ejection fraction | 120
thin rim of pericardial effusion | 120
bilateral moderate pleural effusion | 120
basal atelectasis | 120
discharged from ICU | 168
treated with dexamethasone | 168
improved | 192
generalised oedema subsided | 192
skin rash resolved | 192
conjunctivitis resolved | 192
white blood cell count normalised | 192
renal function improved | 192
inflammatory markers normalised | 192
repeat echocardiography showed trace tricuspid regurgitation | 192
improved right ventricular systolic function | 192
normal size of right atrium and ventricle | 192
normal pulmonary artery systolic pressure | 192
discharged home | 240
tapering dose of prednisolone | 240
follow-up | 336
symptoms resolved | 336
general weakness | 336
fatigue | 336
repeat echocardiogram normal | 336