31 weeks of pregnancy | -672\
emergency cesarean delivery | -672\
abruptio placenta | -672\
birth weight 1090 g | -672\
Apgar values of 4 and 8 in the first and fifth minutes of life | -672\
multiple pregnancy | -672\
hypothyroidism | -672\
gestational diabetes | -672\
group B streptococcal urine infection | -672\
antibiotics | -672\
respiratory distress | 0\
respiration rate of 65 breaths per min | 0\
chest retraction | 0\
CPAP machine | 0\
positive end expiratory pressures | 0\
30% inspired oxygen | 0\
cloudy eyes | 0\
ectropion | 0\
dry ichthyotic skin | 0\
typical male genitalia | 0\
bilaterally undescended testicles | 0\
height 75th percentile | 0\
weight 25th percentile | 0\
head circumference 25th percentile | 0\
temperature 36.2°C | 0\
neurologically fine | 0\
heart rate 167 beats per min | 0\
pulsations well felt | 0\
breath sounds from both sides of the lung equal | 0\
no organomegaly in the abdomen | 0\
normal blood count | 0\
normal electrolytes | 0\
normal liver function | 0\
respiratory distress syndrome | 0\
ground-glass opacity | 0\
minor respiratory acidosis | 0\
surfactant dosage | 12\
CPAP assistance | 12\
bowel movement | 12\
trophic feeding | 72\
breast milk | 72\
abdominal distension | 144\
tachycardia | 144\
tachypnea | 144\
thrombocytopenia | 144\
neutropenia | 144\
raised C-reactive protein level | 144\
meropenem | 144\
vancomycin | 144\
stop the tropic feeding | 216\
negative culture results | 216\
restart feeding | 216\
high-flow oxygen treatment | 336\
relapses of unexplained apnea | 504\
CPAP | 504\
septic examination negative | 504\
normal brain MRI | 504\
nasogastric tube | 504\
occasional breast milk | 504\
preterm formula | 504\
no pale stools | 504\
neonatal cholestasis workup | 504\
conjugated hyperbilirubinemia | 504\
total bilirubin 69.8 umol/L | 504\
negative septic workups | 504\
genetic studies | 504\
progressive familial intrahepatic cholestasis | 504\
ALGS | 504\
normal X-ray of the spine | 504\
normal echocardiogram | 504\
normal eye test | 504\
craniosynostosis | 504\
hepatosplenomegaly not seen | 504\
no signs of biliary atresia | 504\
normal-appearing gallbladder | 504\
no signs of intrahepatic or extrahepatic biliary tree dilatation | 504\
decline in albumin level | 504\
rise in bilirubin | 504\
rise in AST | 504\
rise in ALT | 504\
multiple albumin infusions | 504\
worsening cholestasis | 504\
infectious etiology investigation | 504\
unremarkable results | 504\
normal TSH | 504\
normal T3 | 504\
normal T4 | 504\
normal cortisol | 504\
negative metabolic disorders | 504\
negative galactosemia | 504\
negative tyrosinemia type 1 | 504\
no micropenis | 504\
no hypoglycemia | 504\
whole genomic sequence | 504\
caffeine | 504\
hemoglobin optimization | 504\
phenobarbitone | 504\
severe cyanosis | 936\
apnea | 936\
bradycardia | 936\
aggressive cardio-respiratory resuscitation | 936\
intubation | 936\
mechanical breathing | 936\
epinephrine | 936\
septic shock | 936\
multiorgan failure | 936\
disseminated intravascular coagulation | 936\
acute renal damage | 936\
capillary leak syndrome | 936\
death | 2400\
whole-exome sequencing results | 2400\
pathogenic heterozygous variant c.1076c>T (Ser359Phe) chr1: 120512166 | 2400\
NOTCH2 gene | 2400\
ALGS2 | 2400