57 years old | 0
woman | 0
type 2 diabetes | 0
HbA1c 148 mmol/mol | 0
presented to the emergency department | 0
lower back pain | 0
absence of trauma | 0
right hallux apical neuropathic ulcer | -2928
osteomyelitis | -2928
non-healing wound | -8760
left forefoot amputation | -8760
left fifth toe ulcer | -12528
peripheral vascular disease | 0
peripheral neuropathy | 0
diabetic retinopathy | 0
diabetic nephropathy | 0
atrial fibrillation | 0
hypertension | 0
WHO performance status score 2 | 0
Metformin MR 1 g twice-daily | 0
Lantus 18 units at night | 0
aspirin 75 mg once-daily | 0
bisoprolol 7.5 mg once-daily | 0
cholecalciferol 20 000 units once week | 0
ramipril 5 mg once-daily | 0
rivaroxaban 20 mg once-daily |:0
acutely confused | 0
septic | 0
denied headache | 0
denied respiratory symptoms | 0
denied urinary symptoms | 0
denied gastrointestinal symptoms | 0
BP 102/84 mmHg | 0
heart rate 110/min | 0
temperature 33.7°C | 0
normal heart sounds | 0
no added murmurs | 0
chest clear on auscultation | 0
abdominal examination unremarkable | 0
left foot amputation wound site soft tissue infection | 0
capillary refill time 3 s | 0
biphasic Doppler signals on both posterior tibial arteries | 0
right hallux ulcer dry | 0
no signs of acute infection | 0
lumbar vertebral tenderness | 0
bilateral lower limb weakness | 0
absent reflexes | 0
acute renal failure | 0
profound metabolic acidosis | 0
oliguria | 0
pH 7.13 | 0
pCO2 4.2 kPa | 0
lactate 14.6 mmol/L | 0
bicarbonate 10.3 mmol/L | 0
base excess −18.9 mmol/L | 0
normal chest radiograph | 0
negative urine cultures | 0
CT scan of head no acute intracranial haemorrhage | 0
CT scan of head no collection | 0
CT scan of head no infarct | 0
FAST scan collapsible IVC | 0
FAST scan poorly filled RV | 0
FAST scan excluded abdominal free fluid | 0
FAST scan excluded AAA | 0
CT abdomen no intra-abdominal collections | 0
CT abdomen no source of sepsis | 0
duplex ultrasound diffusely diseased arteries | 0
no haemodynamically significant stenosis in right leg | 0
biphasic spectral waveforms in right lower limb | 0
left leg 50–55% haemodynamically significant stenosis | 0
left mid SFA stenosis | 0
left mid popliteal artery stenosis | 0
crural arteries dense calcification | 0
left lower limb distal anterior tibial artery flow from peroneal artery | 0
triphasic spectral waveforms at left CFA | 0
tri/bi spectral waveforms at left knee | 0
strong monophasic signal below left knee | 0
no acute revascularisation deemed necessary | 0
left forefoot amputation site wound swabs mixed growth | 0
Pseudomonas sp. | 0
yeast | 0
right foot wound swabs negative | 0
previous foot ulcer swabs mixed anaerobes | 0
S. aureus | 0
blood cultures Beta haemolytic group B Streptococcus | 0
transthoracic echocardiogram no vegetations | 0
severely impaired systolic function | 0
EF 25–30% | 0
too unwell for transoesophageal echocardiogram | 0
abdominal imaging unremarkable | 0
spinal MRI arranged | 0
severe sepsis | 0
treated with IV Ceftriaxone | 0
treated with metronidazole | 0
glycaemic control optimized with insulin infusion | 0
vascular team review | 0
concurred with IV antibiotics | 0
no immediate indication for debridement | 0
no immediate indication for surgery | 0
multi-organ failure | 0
severe LVF | 0
acute kidney injury | 0
ischaemic liver dysfunction | 0
MRI confirmed L3/L4 discitis | 0
MRI confirmed L4/L5 discitis | 0
adjacent vertebral end-plate oedema | 0
posterior epidural collection | 0
canal compression extending from T12 to L4 | 0
managed conservatively with antibiotics | 0
ciprofloxacin | 0
gentamicin | 0
meropenem | 0
ceftriaxone | 0
neurosurgical intervention deemed high risk | 0
declined surgery | 0
inflammatory markers improved | 0
remained bed bound | 0
persistent lower limb neurology | 0
further signs of sepsis | 0
passed away | 876
septicaemia | 876
epidural abscess | 876
diabetic foot ulcer | 876
