13 years old | 0
female | 0
admitted to the hospital | 0
fever | -120
productive cough | -120
hemoptysis | -120
diarrhea | -120
alert | 0
respiratory distress | 0
tachycardia | 0
chest indrawing | 0
decreased lung sound on the right side | 0
lymphopenia | 0
elevated C-reactive protein | 0
elevated procalcitonin | 0
elevated lactate dehydrogenase | 0
chest computed tomography scan | 0
nasopharyngeal swab sample collected for RT-PCR test | 0
confirmed diagnosis of COVID-19 | 0
BiPAP | 0
admitted to ICU | 0
Atazanavir | 0
interferon beta-1a | 0
signs worsened | 0
arterial oxygen saturation decreased | 0
plasmapheresis performed four times | 0
fresh-frozen plasma as replacement fluid | 0
elevated WBC count | 0
predominance of PMNs | 168
leukocytosis | 168
chest X-ray revealed significant change in lungs | 48
general condition improved | 48
arterial oxygen saturation improved to 94% | 48
interferon beta-1a injected every 48 hours | 72
tachypnea disappeared | 120
tachycardia disappeared | 120
transferred from ICU to ward | 192
oxygen therapy changed to nasal cannula | 216
respiratory distress disappeared gradually | 216
supplemental oxygen tapered | 216
discharged | 336
normal oxygen saturation in room air | 336
no fever | 336
good condition in 2-week follow-up | 336
platelet count normal | 0
elevated D-Dimer | 0
liver function tests abnormal | 48
bilirubin level abnormal | 48
elevated ferritin | 168
elevated ESR | 168
elevated creatinine | 0
normal pH | 0
normal bicarbonate | 0
normal pCO2 | 0
no problem in follow-up | 336
