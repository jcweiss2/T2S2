74 years old| 0
male| 0
asthma| -87600
nephrotic syndrome| -87600
prednisolone 10 mg daily| -87600
long-term steroid use| -87600
steroid-induced diabetes mellitus| -87600
obesity| -87600
never drank alcohol| 0
never smoked| 0
unconscious state| 0
Glasgow Coma Scale E2V1M4| 0
blood pressure no measurable| 0
carotid artery pulsation present| 0
heart rate 110 beats per minute| 0
respiratory rate 24 breaths per minute| 0
body temperature 35.2°C| 0
body mass index 28| 0
obesity| 0
near obstruction of airway| 0
left conjugated deviated ocular position| 0
right hemiparesis| 0
hematemesis| 0
double incontinence| 0
complete phimosis| 0
hypogonadism| 0
rapid fluid resuscitation| 0
tracheal intubation| 0
mechanical ventilation| 0
nasogastric tube placement| 0
noradrenaline infusion| 0
vasopressin infusion| 0
sinus tachycardia| 0
complete right bundle branch block| 0
atrophic liver| 0
multiple pancreatic cysts| 0
excess visceral fat| 0
penis buried under subcutaneous fat| 0
blood test results available| 0
septic shock of unknown focus| 0
acute respiratory failure| 0
renal failure| 0
hyperkalemia| 0
cerebral ischemia| 0
liver cirrhosis| 0
rhabdomyolysis| 0
diabetes mellitus| 0
upper gastrointestinal bleeding| 0
calcium chloride infusion| 0
insulin therapy| 0
zirconium for hyperkalemia and hyperglycemia| 0
broad-spectrum antibiotics administration| 0
meropenem 2 g per day| 0
linezolid 1200 mg per day| 0
mineral corticoid for septic shock| 0
external urethral orifice unidentified| 0
emergency circumcision| 0
balloon catheter insertion| 0
intensive care unit admission| 0
circulation stabilized| 72
cardiopressor treatment discontinued| 72
PaO2/FiO2 >300| 72
obey orders| 72
extubation| 72
communication with patient| 72
past history confirmed| 72
Staphylococcus capitis blood culture| 72
steroid dose rapidly decreased| 72
circulation became unstable| 72
steroid dose gradually tapered| 72
adrenal insufficiency suspected| 72
ACTH level 5 pg/mL| 72
cortisol level 7.0 μg/dL| 72
adrenal insufficiency confirmed| 72
hepatitis B negative| 72
hepatitis C negative| 72
autoimmune antibodies negative| 72
M2BPGI value 2+| 72
NAFLD fibrosis score 2.0| 72
FIB-4 index 9.45| 72
burn-out NASH diagnosed| 72
ascites| 144
abdominal CT showed ascites| 144
no fresh ischemic lesions| 144
pituitary gland normal appearance| 144
transient ischemic attack| 144
Todd's paralysis| 144
testosterone low| 144
estradiol high| 144
hypogonadism induced by NASH| 144
self-feeding| 168
transfer assistance required| 168
severe lower extremity muscle weakness| 168
disuse| 168
critical illness myopathy| 168
respiratory function deteriorated| 360
enhanced CT showed thrombosis right pulmonary artery| 360
thrombosis right common iliac vein| 360
heparinization| 360
renal function returned to normal| 360
rhabdomyolysis resolved| 360
liver dysfunction| 360
coagulopathy| 360
anemia| 360
left leg phlegmon| 432
antibiotics treatment for phlegmon| 432
esophagogastoscopy showed atrophic gastritis| 648
transferred to another hospital| 816
phlegmon improved| 816
burn-out NASH developed under long-term steroid use| 0
adrenal insufficiency| 72
immune suppression| 0
sepsis with multiple organ failure| 0
pulmonary embolism| 360
gait disturbance due to disuse or critical illness myopathy| 168
leg phlegmon| 432
