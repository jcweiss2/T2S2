53 years old| 0
male| 0
presented to the emergency room| -72
fever| -72
myalgia| -72
confusion| -24
severe frontal headache| -24
no history of sick contacts| 0
no recent travels| 0
no recreational use of drug| 0
no history of chronic alcoholism| 0
no diabetes| 0
no chronic kidney disease| 0
no cardiac disease| 0
no recent throat infection| 0
no skin infection| 0
became more confused and lethargic| 0
lying in bed| 0
moderate distress| 0
Glasgow Coma Scale score of 10| 0
could not follow commands| 0
neck rigidity on flexion| 0
rigidity in the left upper extremity| 0
increased tone on the left side| 0
white blood cell count of 10×10^9/L| 0
hemoglobin level of 13.4 g/dl| 0
thrombocytopenia| 0
platelet count of 54×10^9/L| 0
sodium level of 134 mEq/l| 0
calcium level of 8.4 mg/dl| 0
magnesium level of 1.7 mg/dl| 0
phosphorus level of 3.2 mg/dl| 0
bicarbonate level of 24 mEq/l| 0
blood glucose level of 142 mg/dl| 0
troponin level increased from 0.16 ng/ml–0.38 ng/ml| 0
normal sinus rhythm on ECG| 0
ammonia level of 47 mcmol/l| 0
normal thyroid-stimulating hormone level| 0
normal liver function tests| 0
negative for flu| 0
negative for respiratory syncytial virus| 0
negative for coronavirus disease 2019| 0
negative urine analysis| 0
negative urine toxicology screen| 0
negative salicylate level| 0
negative alcohol level| 0
lumbar puncture performed| 0
elevated white blood cell count of 682×10^9/l| 0
neutrophil 81%| 0
red blood cell count of 10×10^9/l| 0
protein level of 117 mg/dl| 0
glucose level of 58 mg/dl| 0
admitted to the MICU| 0
empirical therapy for meningitis| 0
vancomycin| 0
cefepime 2 g every 8 h| 0
ampicillin 2 g every 4 h| 0
developed new-onset left-sided weakness| 24
computed tomography scan showed no intracranial hemorrhage| 24
incidental finding of 778 mm mass concerning an aneurysm| 24
Methicillin-sensitive staphylococcal aureus in the blood| 24
antibiotics deescalated to Oxacillin 2 g| 24
steroid stopped| 24
transesophageal echo showed vegetation in the aortic valve| 24
intubated for respiratory distress| 24
persistently bacteremic| 24
febrile| 24
ceftaroline added| 24
MRI showed large posterior cerebral artery infarct| 24
consulted cardiothoracic surgery team for aortic valve replacement| 24
surgery not deemed appropriate| 24
repeat computed tomography head scan showed intraparenchymal bleed| 24
lactic acid level rising| 24
worsening kidney function| 24
bicarbonate administered| 24
oxygen saturation levels decreased to 40%| 24
cardiac arrest| 24
cardiopulmonary resuscitation initiated| 24
advanced life support measures employed| 24
pronounced dead| 24
bacterial meningitis secondary to infective endocarditis| 0
Staphylococcus aureus meningitis| 0
infective endocarditis with vegetation| 0
large posterior cerebral artery infarct| 0
intraparenchymal bleed in the right frontal area| 24
embolic stroke| 0
aortic valve vegetation| 0
persistent bacteremia| 24
persistent fever| 24
respiratory distress| 24
acute kidney injury| 24
Methicillin-sensitive Staphylococcal Aureus bacteremia| 24
neurological complications| 0
meningitis| 0
stroke| 0
aortic valve damage| 0
sepsis| 24
death| 24
53 years old|0
male|0
presented to the emergency room|-72
fever|-72
myalgia|-72
confusion|-24
severe frontal headache|-24
no history of sick contacts|0
no recent travels|0
no recreational use of drug|0
no history of chronic alcoholism|0
no diabetes|0
no chronic kidney disease|0
no cardiac disease|0
no recent throat infection|0
no skin infection|0
became more confused and lethargic|0
lying in bed|0
moderate distress|0
Glasgow Coma Scale score of 10|0
could not follow commands|0
neck rigidity on flexion|0
rigidity in the left upper extremity|0
increased tone on the left side|0
white blood cell count of 10×10^9/L|0
hemoglobin level of 13.4 g/dl|0
thrombocytopenia|0
platelet count of 54×10^9/L|0
sodium level of 134 mEq/l|0
calcium level of 8.4 mg/dl|0
magnesium level of 1.7 mg/dl|0
phosphorus level of 3.2 mg/dl|0
bicarbonate level of 24 mEq/l|0
blood glucose level of 142 mg/dl|0
troponin level increased from 0.16 ng/ml–0.38 ng/ml|0
normal sinus rhythm on ECG|0
ammonia level of 47 mcmol/l|0
normal thyroid-stimulating hormone level|0
normal liver function tests|0
negative for flu|0
negative for respiratory syncytial virus|0
negative for coronavirus disease 2019|0
negative urine analysis|0
negative urine toxicology screen|0
negative salicylate level|0
negative alcohol level|0
lumbar puncture performed|0
elevated white blood cell count of 682×10^9/l|0
neutrophil 81%|0
red blood cell count of)10×10^9/l|0
protein level of 117 mg/dl|0
glucose level of 58 mg/dl|0
admitted to the MICU|0
empirical therapy for meningitis|0
vancomycin|0
cefepime 2 g every 8 h|0
ampicillin 2 g every 4 h|0
developed new-onset left-sided weakness|24
computed tomography scan showed no intracranial hemorrhage|24
incidental finding of 778 mm mass concerning an aneurysm|24
Methicillin-sensitive staphylococcal aureus in the blood|24
antibiotics deescalated to Oxacillin 2 g|24
steroid stopped|24
transesophageal echo showed vegetation in the aortic valve|24
intubated for respiratory distress|24
persistently bacteremic|24
febrile|24
ceftaroline added|24
MRI showed large posterior cerebral artery infarct|24
consulted cardiothoracic surgery team for aortic valve replacement|24
surgery not deemed appropriate|24
repeat computed tomography head scan showed intraparenchymal bleed|24
lactic acid level rising|24
worsening kidney function|24
bicarbonate administered|24
oxygen saturation levels decreased to 40%|24
cardiac arrest|24
cardiopulmonary resuscitation initiated|24
advanced life support measures employed|24
pronounced dead|24
bacterial meningitis secondary to infective endocarditis|0
Staphylococcus aureus meningitis|0
infective endocarditis with vegetation|0
large posterior cerebral artery infarct|0
intraparenchymal bleed in the right frontal area|24
embolic stroke|0
aortic valve vegetation|0
persistent bacteremia|24
persistent fever|24
respiratory distress|24
acute kidney injury|24
Methicillin-sensitive Staphylococcal Aureus bacteremia|24
neurological complications|0
meningitis|0
stroke|0
aortic valve damage|0
sepsis|24
death|24
