17 years old | 0
male | 0
complete transposition of the great arteries | -7200
ventricular septal defect | -7200
pulmonary stenosis | -7200
Rastelli repair | -7200
placement of a 16 mm pulmonary homograft | -7200
conduit replacement with a 20 mm aortic homograft | -5040
balloon dilated | -2160
transcatheter Melody valve placement | -2160
fever | -48
diarrhea | -48
vomiting | -48
syncope | -48
admitted to the intensive care unit | 0
pale | 0
febrile | 0
icteric | 0
tachycardic | 0
hypotensive | 0
blood cultures grew methicillin-sensitive staphylococcus aureus | 0
intravenous fluids | 0
inotropes (dopamine 5 μg/kg/min) | 0
intravenous vancomycin (1 g every 12 h) | 0
rifampicin (300 mg every 8 h) | 0
gentamicin (62 mg every 12 h) | 0
vancomycin stopped | 12
intravenous oxacillin (2 g every 4th h) | 12
right ventricular pressure estimates on echocardiography were initially normal | 0
increased right ventricular pressure estimates on echocardiography | 24
cardiac magnetic resonance (CMR) imaging | 24
computed tomography (CT) of the chest | 24
multiple cavitary nodules of varying sizes throughout both the lungs | 24
septic emboli | 24
condition stabilized | 48
discharged from the intensive care unit | 48
gentamicin stopped | 336
explantation of the Melody valve | 432
inflammation around the heavily calcified homograft | 432
Melody valve was clearly infected | 432
thickening and edema of both the valve leaflets | 432
valve leaflets adhered to the internal wall of the Melody valve | 432
homograft and Melody valve explanted | 432
replaced with a pulmonary homograft | 432
histopathological examination revealed acute inflammatory infiltrate | 432
granulation tissue in the Melody valve | 432
postoperative course was uneventful | 432
doing well at 6 months follow-up | 2160