22 years old | 0
male | 0
admitted to the hospital | 0
5-year history of smoking | -8760
exposed to live poultry | -48
high fever | -72
chills | -72
ibuprofen | -72
azithromycin | -72
visit to the local hospital | -72
complaints progressed | -48
visit to the emergency department | 0
lymphopenia | 0
thrombocytopenia | 0
normal white blood cell count | 0
normal PaO2/FiO2 values | 0
patchy shadows and consolidation in the lower lobe of the right lung | 0
meropenem | 0
moxifloxacin | 0
throat swab sample obtained | -24
oseltamivir | -24
PaO2/FiO2 value declined | 24
septic shock | 24
SOFA score increased | 24
H5N6 virus identified | 24
transferred to the ICU | 24
invasive mechanical ventilation | 24
low tidal volume | 24
open lung ventilation strategy | 24
bronchoalveolar lavage fluid galactomannan test | 24
dosage of oseltamivir increased | 24
peramivir | 24
amphotericin B | 24
low-dose corticosteroid | 24
mediastinal and subcutaneous emphysema | 120
CT images showed rapid progression of lung consolidation | 168
venovenous extracorporeal membrane oxygenation | 168
sirolimus | 192
viral titer of the tracheal aspirate sample | 192
viral titers decreased | 216
H5N6 virus undetectable in throat swab specimens | 240
H5N6 virus undetectable in tracheal aspirate samples | 312
ECMO stopped | 336
endotracheal tube removed | 336
sirolimus, NAIs, and antibiotics discontinued | 336
discharged | 468
follow-up | 1752
bilateral interstitial changes in the lungs | 1752
pulmonary function test showed normal ventilation | 1752
slightly decreased efficiency in diffusion | 1752