66 years old | 0
male | 0
Type II diabetes mellitus | 0
hypertension | 0
hyperlipidemia | 0
admitted to the hospital | 0
acute shortness of breath | -24
cough | -24
fever | -24
travel history to Batam, Indonesia | -24
temperature 38.0°C | 0
blood pressure 130/70 mmHg | 0
pulse 140 bpm | 0
respiratory rate of 25 per minute | 0
oxygen saturation 92% on room air | 0
placed on a 40% Venturi mask | 0
bilateral crepitations | 0
20 × 20 cm back carbuncle | 0
white blood cell count of 31000/µl | 0
hemoglobin level of 11. 5 g/dl | 0
lactate level of 5.92 mmol/L | 0
pro-brain natriuretic peptide level of 731 pg/ml | 0
arterial blood gas in supplemental oxygen showed a pH level of 7.42 | 0
pCO2 of 35.1 mmHg | 0
pO2 of 91.9 mmHg | 0
PaO2/FiO2 ratio of 230 | 0
chest X-ray (CXR) revealed bilateral diffuse pulmonary infiltrates | 0
saucerization of the carbuncle | 0
surgery | 0
COVID-19 swab test | 0
team huddle | 0
transportation of the patient to the operating theatre (OT) | 0
signages posted | 0
security personnel deployed | 0
plastic cover on the trolley removed and discarded into a biohazard bag | 0
airway trolley placed in the OT | 0
C-Mac video laryngoscope with disposable blade | 0
preoxygenation | 0
modified rapid sequence induction | 0
induction agents administered | 0
mask ventilation avoided | 0
intubation | 0
general anesthesia maintained with desflurane | 0
mechanical ventilation with a tidal volume of 7 ml/kg | 0
patient kept intubated | 0
COVID-19 test result negative | 24
discharged | 24