32 years old|0
man|0
presented at the Emergency Department|0
tonic-clonic seizures|0
hypoxemia|0
admitted to the Intensive Care Unit|0
endotracheal tube placed|0
invasive mechanical ventilation initiated|0
sedation with midazolam|0
fentanyl for analgesia|0
chest X-ray showed right basal atelectatic band|0
computed tomography (CT) scan of the chest showed bilateral basal condensation areas|0
brain CT scan showed normal brain|0
hypothyroidism|0
levothyroxine|0
morbid type 3 obesity|0
gastritis|0
gastric ulcer|0
penicillin allergies|0
endoscopic procedure for erosive gastropathy|-168
piperacillin plus tazobactam initiated|0
clindamycin initiated|0
sputum samples taken for cultures|0
blood samples taken for cultures|0
urine samples taken for cultures|0
day 2 in the ICU|48
remained sedated with midazolam|48
fentanyl for analgesia continued|48
day 3 in the ICU|72
bronchoscopy performed|72
reddened mucosa with cavity|72
hemorrhagic stitches|72
active bleeding|72
bronchioalveolar lavage samples analyzed|72
MRSA identified|72
mecA gene-resistance mechanism|72
luk-PV gene-resistance mechanism|72
piperacillin plus tazobactam suspended|72
intravenous vancomycin administered|72
cerebrospinal fluid obtained by lumbar puncture|0
no bacterial growth in cerebrospinal fluid|0
day 4 in the ICU|96
significant clinical improvement|96
weaning of sedation initiated|96
weaning of invasive mechanical ventilation initiated|96
extubated|96
good ventilatory mechanics|96
99% saturation|96
oxygen support with mask initiated|96
respiratory rate of 19 breaths/min|96
oriented to time, space, and person|96
Glasgow Coma Scale score of 15/15|96
reactive isochoric pupils|96
day 5 in the ICU|120
afebrile|120
awake|120
breathing ambient air|120
day 6 in the ICU|144
discharged from ICU|144
remained hospitalized|144
discharged after 10-day hospital stay|240
followed up in Outpatient Department|240
remains in general good health after 6 months|2400
cavitary pneumonia due to MRSA|0
no previous respiratory symptoms|0
no history of tobacco use|0
no illicit drug use|0
no human immunodeficiency virus|0
no nasopharyngeal colonization for Staphylococcus|0
no adverse events related to endoscopic procedure|-168
no hospital admission prior to endoscopic procedure|-168
no MRSA infections prior|0
no recent hospitalization|0
no residence in nursing homes|0
no long-term care facilities|0
no medical devices|0
no permanent catheters|0
leukocytes 17 900/mm3|0
neutrophils 85.6%|0
hematocrit 34.3%|0
hemoglobin 11.4 g/dL|0
platelets 280 000/mm3|0
sodium 141.0 mEq/L|0
potassium 3.9 mEq/L|0
chloride 109 mEq/L|0
glucose 125.40 mg/dL|0
blood urea nitrogen 14 mg/dL|0
creatinine 0.7 mg/dL|0
prothrombin time 13.1 s|0
partial thromboplastin time 30.6 s|0
cavitary area in bronchoscopic image|72
hemorrhagic stitches in bronchoscopic image|72
active bleeding area in bronchoscopic image|72
response to vancomycin|72
