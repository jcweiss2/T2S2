34 years old | 0
African-American | 0
female | 0
admitted to the hospital | 0
menorrhagia | -672
pelvic pain | -672
left uterine mass | -672
myoma | -672
ultrasound | -672
multiple small myomas | -672
diagnostic laparoscopy | 0
myomectomy | 0
past surgical history | -10080
laparotomy | -10080
left oophorectomy | -10080
ovarian cysts | -10080
elective terminations of pregnancy | -10080
inflammatory process | -10080
asthma | -10080
nonsteroidal anti-inflammatory drugs | -10080
physical examination | 0
bradycardia | 0
thyroid nodule | 0
laboratory workup | 0
mild iron deficiency anemia | 0
inconclusive thyroid studies | 0
euthyroid | 0
open entry method | 0
adherent small bowel loops | 0
pneumoperitoneum | 0
exploration of the abdomen | 0
extensive adhesions | 0
port placement | 0
adhesiolysis | 0
disposable scissors | 0
pelvic organs | 0
uterus | 0
sigmoid colon | 0
myolysis | 0
bipolar needle punctures | 0
abdomen lavaged | 0
saline | 0
operative time | 0
anesthetic inhalation agents | 0
sevoflurane | 0
nitrous oxide | 0
estimated blood loss | 0
discharged | 0
postoperative recovery | 0
afebrile | 24
voiding well | 24
oral intake | 24
passed flatus | 48
bowel movement | 72
bloody drainage | 24
hydroflation | 24
black and blue mark | 48
abdominal pain | 24
distention | 24
vomited | 96
emergency room | 96
acute abdomen | 96
surgical team | 96
atrial fibrillation | 96
hypotension | 96
triple lumen catheter | 96
operating room | 96
exploratory laparotomy | 96
enteric fluid | 96
umbilical port site | 96
midline laparotomy | 96
gross spillage | 96
adhesions | 96
bowel | 96
anterior abdominal wall | 96
mobilization | 96
small bowel | 96
perforated bowel | 96
enterotomy | 96
adhesiolysis | 96
resected bowel | 96
Prasad double barrel ileostomy | 96
pathology report | 96
ischemic necrosis | 96
bowel mucosa | 96
edematous | 96
intensive care unit | 96
broad-spectrum antibiotics | 96
activated protein C | 96
Xigris | 96
candidemia | 120
unsuccessful extubation trials | 120
multiple neuropathy | 120
nosocomial pneumonia | 120
pressure ulcer | 120
drug-induced thrombocytopenia | 120
gastrointestinal bleeding | 120
shock | 120
cardiopulmonary arrests | 120
gastrostomy | 120
tracheostomy | 120
inferior vena cava filter | 120
deep-vein thrombosis | 120
rehabilitation | 744