63 years old | 0
male | 0
admitted to the hospital | 0
feeling unwell | -336
vancomycin resistant enterococcal | 0
dehiscence of the aortic valve | 0
aortic valve root abscess | 0
mitral valve vegetations | 0
patent foramen ovale | 0
inferior vena cava Eustachian valve | 0
liver failure | 0
renal failure | 0
bilirubin 54 mg/dL | 0
alkaline phosphatase 222 IU/L | 0
alanine aminotransferase 1211 IU/L | 0
continuous veno-venous hemofiltration | 0
heparin as anticoagulant | 0
platelet count 179 × 10^3 per mm^3 | 0
drop in platelet count to 35 × 10^3 per mm^3 | 72
heparin induced thrombocytopenia | 72
heparin stopped | 72
Danaparoid as hemofiltration anticoagulation | 72
platelet counts dropped to 16 × 10^3 per mm^3 | 168
aortic valve replacement | -672
Aspirin | -672
bisoprolol | -672
perindopril | -672
atorvastatin | -672
redo-aortic valve replacement | 0
mitral valve repair | 0
closure of the patent foramen ovale | 0
repair of the aortic root abscess | 0
excision of the Eustachian valve | 0
ventilator dependence | 0
tracheostomy | 0
renal replacement therapy | 0
cardiovascular support | 0
milrinone 10 ml/h | 0
noradrenaline 20 ml/h | 0
vasopressin 2 IU/h | 0
discharged | 4320
SDF device used | 48
sub-lingual microvasculature examined | 48
sepsis | 48
pyrexia | 48
low systemic vascular resistance | 48
increased inflammatory markers | 48
increased inotropic-vasoconstrictor support | 48
HIT | 48
vessel density measured | 48
perfusion quality measured | 48
TVD 20.35 | 48
PVD 17.25 | 48
De Backer score 11.66 | 48
PPV 83.69 | 48
MFI 1 | 48
FHI 0 | 48
CI 3.7 | 48
MAP 66 | 48
SVRI 1038 | 48
pH 7.42 | 48
lactate 4.9 | 48
noradrenaline 0.3 | 48
vasopressin 1 | 48
SDF device used | 60
sub-lingual microvasculature examined | 60
vessel density measured | 60
perfusion quality measured | 60
TVD 37.21 | 60
PVD 37.21 | 60
De Backer score 21.37 | 60
PPV 100 | 60
MFI 3.5 | 60
FHI 0.28 | 60
CI 2.9 | 60
MAP 55 | 60
SVRI 1178 | 60
pH 7.36 | 60
lactate 6.9 | 60
noradrenaline 0.2 | 60
vasopressin 1 | 60
SDF device used | 90
sub-lingual microvasculature examined | 90
vessel density measured | 90
perfusion quality measured | 90
TVD 35.78 | 90
PVD 35.78 | 90
De Backer score 22.54 | 90
PPV 100 | 90
MFI 3 | 90
FHI 0 | 90
CI 2.8 | 90
MAP 74 | 90
SVRI 1885 | 90
pH 7.2 | 90
lactate 6.6 | 90
noradrenaline 0.26 | 90
vasopressin 4 | 90
SDF device used | 1104
sub-lingual microvasculature examined | 1104
vessel density measured | 1104
perfusion quality measured | 1104
TVD 36.86 | 1104
PVD 36.86 | 1104
De Backer score 22.39 | 1104
PPV 100 | 1104
MFI 3 | 1104
FHI 0 | 1104
CI 2.8 | 1104
MAP 52 | 1104
SVRI 1715 | 1104
pH 7.45 | 1104
lactate 1.1 | 1104
noradrenaline 0.06 | 1104
vasopressin 0 | 1104