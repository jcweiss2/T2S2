66 years old | 0
female | 0
admitted to the hospital | 0
mild cough | -48
sore throat | -48
asthma | -672
fever | -24
dialysis session | -24
COVID-19 positive | 0
droplet and contact isolation precautions | 0
productive cough | 0
dyspnea | 12
oxygen saturation 86% | 12
oxygen 2 L/min by nasal cannula | 12
respiratory deterioration | 24
intubated | 24
septic shock | 24
ceftriaxone | 24
ciprofloxacin | 24
hydroxychloroquine | 24
NP swab negative for influenza | 24
oseltamivir not treated | 24
continuous renal replacement therapy (CRRT) | 48
regional citrate anticoagulation | 48
critical care nursing staff training | 48
care bundle approach | 48
CRRT dosing reduced | 48
extubated | 456
discharged home | 480
readmitted | 888
biliary obstruction | 888
biochemistry | 888
endoscopic retrograde cholangiopancreatographies | 888
critical illness-associated secondary sclerosing cholangitis | 888
infected liver abscesses | 888
antimicrobial therapy | 888
fluconazole | 888
moxifloxacin | 888
contact tracing | 24
staff exposed | 24
HD patients exposed | 24
self-isolation | 24
surveillance NP swabs | 24
negative NP swabs | 24
cleared to return to work | 168
universal PPE precautions | 744
mask and visor | 744
asymptomatic staff members | 744
no self-isolation | 744
essential visitors screened | 744
mask required | 744
dialysis patients informed | 744
printed letter | 744
updated signs | 744
PDSA cycles | 744
COVID-19 screening evolution | 744
infectious disease specialists | 744
infection control practitioners | 744
local disease transmission patterns | 744
COVID-19 Nephrology task force | 744
daily review | 744
IP & C | 744
hospital-wide policy | 744
Canadian Society of Nephrology COVID-19 Rapid Response Team | 744
national information | 744
international collaboration | 744
Wang et al | 744
HD patients with COVID-19 | 744
nonrespiratory complaints | 744
abdominal pain | 744
diarrhea | 744
screening protocols | 744
model for improvement framework | 744
rapid PDSA cycles | 744
evolving information | 744
disease symptoms | 744
spread | 744
future screening protocols | 744
lessons learned | 744
vulnerable populations | 744
in-center HD | 744
quality improvement methodology | 744
rapid PDSA cycles | 744
new knowledge | 744
best practices | 744
limit risks | 744
potential outbreak | 744
dialysis unit | 744
acute complications | 744
delayed complications | 744
COVID-19 | 744