29 years old | 0
male | 0
admitted to the hospital | 0
deafness | -103008
severe headaches | -72
confusion | -72
visual disorders | -72
temporospatial disorientation | 0
incomplete ophthalmologic examination | 0
scheduled fundoscopic examination with retinal fluorescein angiography | 0
perception hearing disorder | -103008
bilateral sensorineural deafness | 0
slight elevated protein level in CSF | 0
lymphocytic pleocytosis in CSF | 0
normal glucose level in CSF | 0
negative oligoclonal bands in CSF | 0
unremarkable laboratory tests | 0
negative blood screening for infections and vasculitis | 0
normal angio-CT | 0
brain MRI with multiple small lesions in corpus callosum | 0
periventricular lesions in hemispheres | 0
deep gray nuclei lesions | 0
midbrain lesions | 0
high-signal abnormalities on T2 and FLAIR sequences | 0
no restriction on DWI | 0
no enhancement on T1 post-contrast | 0
evoked Susac syndrome | 0
neurological status worsened | 0
second MRI showing extensive lesions | 168
instituted corticosteroid therapy (methylprednisolone) | 0
intravenous immunoglobulin pulse | 0
became unconscious | 168
respiratory distress | 168
transfer to intensive care | 168
intubated | 168
complicated by sepsis | 168
limited use of immunosuppressive drugs | 168
death | 1680
