54 years old | 0
female | 0
farmer | 0
admitted to the hospital | 0
7-day history of fever | -168
myalgia | -168
fatigue | -168
poor oral intake | -168
climbed a mountain | -336
treated with antipyretics | -168
fluid therapy | -168
symptoms not relieved | -120
became somnolent | -96
could not follow commands | -96
thrombocytopenia | -96
leukopenia | -96
elevated aspartate aminotransferase | -96
elevated alanine aminotransferase | -96
transferred to hospital | -96
temperature 37.2°C | 0
blood pressure 125/81 mm/Hg | 0
pulse 105 beats per minute | 0
respiratory rate 22 breaths per minute | 0
oxygen saturation 92% | 0
acutely ill | 0
confused | 0
Glasgow coma scale 13 | 0
pupil light reflex normal | 0
no meningeal irritation signs | 0
conjunctivae clear | 0
no palpable lymph nodes | 0
no insect bite site | 0
no eschar | 0
no skin rash | 0
no ecchymosis | 0
mild leucopenia | 0
thrombocytopenia | 0
azotemia | 0
hyperkalemia | 0
elevated liver enzymes | 0
substantially increased creatinine kinase | 0
myoglobin | 0
aldolase | 0
rhabdomyolysis | 0
blood cultures for bacteria negative | 0
serum serology tests negative | 0
reverse transcriptase polymerase chain reaction assay for SFTS virus | 0
plain chest radiograph showed mild pulmonary congestion | 0
bilateral pleural effusion | 0
computed tomography scan of abdomino-pelvis normal | 0
brain CT and magnetic resonance imaging normal | 0
intravenous piperacillin/tazobactam | 0
levofloxacin | 0
emergent continuous renal replacement therapy | 0
metabolic acidosis | 0
hyperkalemia | 0
died | 72
SFTS virus demonstrated | 72
acute respiratory distress syndrome | 72
multiple organ failure | 72
seizure | -96
meningitis | -96
encephalitis | -96
spontaneous intracranial hemorrhage | -96
gadolinium-enhanced brain MRI | 0
lumbar puncture planned | 0
electroencephalography planned | 0
neuromuscular blocker used | 24
muscle enzymes increased | 24
SFTS | 0
myalgia | -168
elevated creatinine kinase | -168
rhabdomyolysis associated with SFTS | 0
influenza | 0
parainfluenza | 0
coxsackievirus | 0
enterovirus | 0
adenovirus | 0
herpes simplex virus | 0
myotoxic cytokines | 0
muscular damage | 0
excessive cytokine production | 0
tissue degeneration | 0
necrosis | 0
regeneration | 0
inflammatory cells | 0
histologic examination | 0
muscle biopsies | 0
SFTS virus | 0
severe disease | 0
overwhelming cytokine production | 0
myalgia | -168
severe myalgia | 0
elevated creatine kinase levels | 0
rhabdomyolysis | 0
SFTS patients | 0
acute febrile diseases | 0
leptospirosis | 0
human granulocytic anaplasmosis | 0
scrub typhus | 0
hemorrhagic fever renal syndrome | 0
co-infection | 0
seizure-like motion | 0
electrolyte disorder | 0
trauma | 0
non-traumatic origin | 0
drug | 0
toxin | 0
seizure | 0
meningitis | 0
encephalitis | 0
spontaneous intracranial hemorrhage | 0
thrombocytopenia | -96
encephalitis or hemorrhage | 0
lumbar puncture | 0
electroencephalography | 0
prone position | 48
rapidly progressive acute respiratory distress syndrome | 48
multiple organ failure | 72
SFTS virus | 72
reverse transcriptase polymerase chain reaction | 72
Korea Centers for Disease Control and Prevention | 72
SFTS case reported in Korea | -876
SFTS cases reported | -876
farmers or forest workers | -876
rural areas | -876
myalgia | -168
fever | -168
thrombocytopenia | -168
month of August | -168
SFTS | 0
rhabdomyolysis | 0
acute febrile diseases | 0
leptospirosis | 0
human granulocytic anaplasmosis | 0
scrub typhus | 0
hemorrhagic fever renal syndrome | 0
co-infection | 0
seizure | -96
meningitis | -96
encephalitis | -96
spontaneous intracranial hemorrhage | -96
thrombocytopenia | -96
encephalitis or hemorrhage | 0
lumbar puncture | 0
electroencephalography | 0
prone position | 48
rapidly progressive acute respiratory distress syndrome | 48
multiple organ failure | 72
SFTS virus | 72
reverse transcriptase polymerase chain reaction | 72
Korea Centers for Disease Control and Prevention | 72
SFTS case reported in Korea | -876
SFTS cases reported | -876
farmers or forest workers | -876
rural areas | -876
myalgia | -168
fever | -168
thrombocytopenia | -168
month of August | -168
SFTS | 0
rhabdomyolysis | 0
acute febrile diseases | 0
leptospirosis | 0
human granulocytic anaplasmosis | 0
scrub typhus | 0
hemorrhagic fever renal syndrome | 0
co-infection | 0
seizure | -96
meningitis | -96
encephalitis | -96
spontaneous intracranial hemorrhage | -96
thrombocytopenia | -96
encephalitis or hemorrhage | 0
lumbar puncture | 0
electroencephalography | 0
prone position | 48
rapidly progressive acute respiratory distress syndrome | 48
multiple organ failure | 72
SFTS virus | 72
reverse transcriptase polymerase chain reaction | 72
Korea Centers for Disease Control and Prevention | 72
SFTS case reported in Korea | -876
SFTS cases reported | -876
farmers or forest workers | -876
rural areas | -876
myalgia | -168
fever | -168
thrombocytopenia | -168
month of August | -168
SFTS | 0
rhabdomyolysis | 0
acute febrile diseases | 0
leptospirosis | 0
human granulocytic anaplasmosis | 0
scrub typhus | 0
hemorrhagic fever renal syndrome | 0
co-infection | 0
seizure | -96
meningitis | -96
encephalitis | -96
spontaneous intracranial hemorrhage | -96
thrombocytopenia | -96
encephalitis or hemorrhage | 0
lumbar puncture | 0
electroencephalography | 0
prone position | 48
rapidly progressive acute respiratory distress syndrome | 48
multiple organ failure | 72
SFTS virus | 72
reverse transcriptase polymerase chain reaction | 72
Korea Centers for Disease Control and Prevention | 72
SFTS case reported in Korea | -876
SFTS cases reported | -876
farmers or forest workers | -876
rural areas | -876
myalgia | -168
fever | -168
thrombocytopenia | -168
month of August | -168
SFTS | 0
rhabdomyolysis | 0
acute febrile diseases | 0
leptospirosis | 0
human granulocytic anaplasmosis | 0
scrub typhus | 0
hemorrhagic fever renal syndrome | 0
co-infection | 0
seizure | -96
meningitis | -96
encephalitis | -96
spontaneous intracranial hemorrhage | -96
thrombocytopenia | -96
encephalitis or hemorrhage | 0
lumbar puncture | 0
electroencephalography | 0
prone position | 48
rapidly progressive acute respiratory distress syndrome | 48
multiple organ failure | 72
SFTS virus | 72
reverse transcriptase polymerase chain reaction | 72
Korea Centers for Disease Control and Prevention | 72
SFTS case reported in Korea | -876
SFTS cases reported | -876
farmers or forest workers | -876
rural areas | -876
myalgia | -168
fever | -168
thrombocytopenia | -168
month of August | -168
SFTS | 0
rhabdomyolysis | 0
acute febrile diseases | 0
leptospirosis | 0
human granulocytic anaplasmosis | 0
scrub typhus | 0
hemorrhagic fever renal syndrome | 0
co-infection | 0
seizure | -96
meningitis | -96
encephalitis | -96
spontaneous intracranial hemorrhage | -96
thrombocytopenia | -96
encephalitis or hemorrhage | 0
lumbar puncture | 0
electroencephalography | 0
prone position | 48
rapidly progressive acute respiratory distress syndrome | 48
multiple organ failure | 72
SFTS virus | 72
reverse transcriptase polymerase chain reaction | 72
Korea Centers for Disease Control and Prevention | 72
SFTS case reported in Korea | -876
SFTS cases reported | -876
farmers or forest workers | -876
rural areas | -876
myalgia | -168
fever | -168
thrombocytopenia | -168
month of August | -168
SFTS | 0
rhabdomyolysis | 0
acute febrile diseases | 0
leptospirosis | 0
human granulocytic anaplasmosis | 0
scrub typhus | 0
hemorrhagic fever renal syndrome | 0
co-infection | 0
seizure | -96
meningitis | -96
encephalitis | -96
spontaneous intracranial hemorrhage | -96
thrombocytopenia | -96
encephalitis or hemorrhage | 0
lumbar puncture | 0
electroencephalography | 0
prone position | 48
rapidly progressive acute respiratory distress syndrome | 48
multiple organ failure | 72
SFTS virus | 72
reverse transcriptase polymerase chain reaction | 72
Korea Centers for Disease Control and Prevention | 72
SFTS case reported in Korea | -876
SFTS cases reported | -876
farmers or forest workers | -876
rural areas | -876
myalgia | -168
fever | -168
thrombocytopenia | -168
month of August | -168
SFTS | 0
rhabdomyolysis | 0
acute febrile diseases | 0
leptospirosis | 0
human granulocytic anaplasmosis | 0
scrub typhus | 0
hemorrhagic fever renal syndrome | 0
co-infection | 0
seizure | -96
meningitis | -96
encephalitis | -96
spontaneous intracranial hemorrhage | -96
thrombocytopenia | -96
encephalitis or hemorrhage | 0
lumbar puncture | 0
electroencephalography | 0
prone position | 48
rapidly progressive acute respiratory distress syndrome | 48
multiple organ failure | 72
SFTS virus | 72
reverse transcriptase polymerase chain reaction | 72
Korea Centers for Disease Control and Prevention | 72
SFTS case reported in Korea | -876
SFTS cases reported | -876
farmers or forest workers | -876
rural areas | -876
myalgia | -168
fever | -168
thrombocytopenia | -168
month of August | -168
SFTS | 0
rhabdomyolysis | 0
acute febrile diseases | 0
leptospirosis | 0
human granulocytic anaplasmosis | 0
scrub typhus | 0
hemorrhagic fever renal syndrome | 0
co-infection | 0
seizure | -96
meningitis | -96
encephalitis | -96
spontaneous intracranial hemorrhage | -96
thrombocytopenia | -96
encephalitis or hemorrhage | 0
lumbar puncture | 0
electroencephalography | 0
prone position | 48
rapidly progressive acute respiratory distress syndrome | 48
multiple organ failure | 72
SFTS virus | 72
reverse transcriptase polymerase chain reaction | 72
Korea Centers for Disease Control and Prevention | 72
SFTS case reported in Korea | -876
SFTS cases reported | -876
farmers or forest workers | -876
rural areas | -876
myalgia | -168
fever | -168
thrombocytopenia | -168
month of August | -168
SFTS | 0
rhabdomyolysis | 0
acute febrile diseases | 0
leptospirosis | 0
human granulocytic anaplasmosis | 0
scrub typhus | 0
hemorrhagic fever renal syndrome | 0
co-infection | 0
seizure | -96
meningitis | -96
encephalitis | -96
spontaneous intracranial hemorrhage | -96
thrombocytopenia | -96
encephalitis or hemorrhage | 0
lumbar puncture | 0
electroencephalography | 0
prone position | 48
rapidly progressive acute respiratory distress syndrome | 48
multiple organ failure | 72
SFTS virus | 72
reverse transcriptase polymerase chain reaction | 72
Korea Centers for Disease Control and Prevention | 72
SFTS case reported in Korea | -876
SFTS cases reported | -876
farmers or forest workers | -876
rural areas | -876
myalgia | -168
fever | -168
thrombocytopenia | -168
month of August | -168
SFTS | 0
rhabdomyolysis | 0
acute febrile diseases | 0
leptospirosis | 0
human granulocytic anaplasmosis | 0
scrub typhus | 0
hemorrhagic fever renal syndrome | 0
co-infection | 0
seizure | -96
meningitis | -96
encephalitis | -96
spontaneous intracranial hemorrhage | -96
thrombocytopenia | -96
encephalitis or hemorrhage | 0
lumbar puncture | 0
electroencephalography | 0
prone position | 48
rapidly progressive acute respiratory distress syndrome | 48
multiple organ failure | 72
SFTS virus | 72
reverse transcriptase polymerase chain reaction | 72
Korea Centers for Disease Control and Prevention | 72
SFTS case reported in Korea | -876
SFTS cases reported | -876
farmers or forest workers | -876
rural areas | -876
myalgia | -168
fever | -168
thrombocytopenia | -168
month of August | -168
SFTS | 0
rhabdomyolysis | 0
acute febrile diseases | 0
leptospirosis | 0
human granulocytic anaplasmosis | 0
scrub typhus | 0
hemorrhagic fever renal syndrome | 0
co-infection | 0
seizure | -96
meningitis | -96
encephalitis | -96
spontaneous intracranial hemorrhage | -96
thrombocytopenia | -96
encephalitis or hemorrhage | 0
lumbar puncture | 0
electroencephalography | 0
prone position | 48
rapidly progressive acute respiratory distress syndrome | 48
multiple organ failure | 72
SFTS virus | 72
reverse transcriptase polymerase chain reaction | 72
Korea Centers for Disease Control and Prevention | 72
SFTS case reported in Korea | -876
SFTS cases reported | -876
farmers or forest workers | -876
rural areas | -876
myalgia | -168
fever | -168
thrombocytopenia | -168
month of August | -168
SFTS | 0
rhabdomyolysis | 0
acute febrile diseases | 0
leptospirosis | 0
human granulocytic anaplasmosis | 0
scrub typhus | 0
hemorrhagic fever renal syndrome | 0
co-infection | 0
seizure | -96
meningitis | -96
encephalitis | -96
spontaneous intracranial hemorrhage | -96
thrombocytopenia | -96
encephalitis or hemorrhage | 0
lumbar puncture | 0
electroencephalography | 0
prone position | 48
rapidly progressive acute respiratory distress syndrome | 48
multiple organ failure | 72
SFTS virus | 72
reverse transcriptase polymerase chain reaction | 72
Korea Centers for Disease Control and Prevention | 72
SFTS case reported in Korea | -876
SFTS cases reported | -876
farmers or forest workers | -876
rural areas | -876
myalgia | -168
fever | -168
thrombocytopenia | -168
month of August | -168
SFTS | 0
rhabdomyolysis | 0
acute febrile diseases | 0
leptospirosis | 0
human granulocytic anaplasmosis | 0
scrub typhus | 0
hemorrhagic fever renal syndrome | 0
co-infection | 0
seizure | -96
meningitis | -96
encephalitis | -96
spontaneous intracranial hemorrhage | -96
thrombocytopenia | -96
encephalitis or hemorrhage | 0
lumbar puncture | 0
electroencephalography | 0
prone position | 48
rapidly progressive acute respiratory distress syndrome | 48
multiple organ failure | 72
SFTS virus | 72
reverse transcriptase polymerase chain reaction | 72
Korea Centers for Disease Control and Prevention | 72
SFTS case reported in Korea | -876
SFTS cases reported | -876
farmers or forest workers | -876
rural areas | -876
myalgia | -168
fever | -168
thrombocytopenia | -168
month of August | -168
SFTS | 0
rhabdomyolysis | 0
acute febrile diseases | 0
leptospirosis | 0
human granulocytic anaplasmosis | 0
scrub typhus | 0
hemorrhagic fever renal syndrome | 0
co-infection | 0
seizure | -96
meningitis | -96
encephalitis | -96
spontaneous intracranial hemorrhage | -96
thrombocytopenia | -96
encephalitis or hemorrhage | 0
lumbar puncture | 0
electroencephalography | 0
prone position | 48
rapidly progressive acute respiratory distress syndrome | 48
multiple organ failure | 72
SFTS virus | 72
reverse transcriptase polymerase chain reaction | 72
Korea Centers for Disease Control and Prevention | 72
SFTS case reported in Korea | -876
SFTS cases reported | -876
farmers or forest workers | -876
rural areas | -876
myalgia | -168
fever | -168
thrombocytopenia | -168
month of August | -168
SFTS | 0
rhabdomyolysis | 0
acute febrile diseases | 0
leptospirosis | 0
human granulocytic anaplasmosis | 0
scrub typhus | 0
hemorrhagic fever renal syndrome | 0
co-infection | 0
seizure | -96
meningitis | -96
encephalitis | -96
spontaneous intracranial hemorrhage | -96
thrombocytopenia | -96
encephalitis or hemorrhage | 0
lumbar puncture | 0
electroencephalography | 0
prone position | 48
rapidly progressive acute respiratory distress syndrome | 48
multiple organ failure | 72
SFTS virus | 72
reverse transcriptase polymerase chain reaction | 72
Korea Centers for Disease Control and Prevention | 72
SFTS case reported in Korea | -876
SFTS cases reported | -876
farmers or forest workers | -876
rural areas | -876
myalgia | -168
fever | -168
thrombocytopenia | -168
month of August | -168
SFTS | 0
rhabdomyolysis | 0
acute febrile diseases | 0
leptospirosis | 0
human granulocytic anaplasmosis | 0
scrub typhus | 0
hemorrhagic fever renal syndrome | 0
co-infection | 0
seizure | -96
meningitis | -96
encephalitis | -96
spontaneous intracranial hemorrhage | -96
thrombocytopenia | -96
encephalitis or hemorrhage | 0
lumbar puncture | 0
electroencephalography | 0
prone position | 48
rapidly progressive acute respiratory distress syndrome | 48
multiple organ failure | 72
SFTS virus | 72
reverse transcriptase polymerase chain reaction | 72
Korea Centers for Disease Control and Prevention | 72
SFTS case reported in Korea | -876
SFTS cases reported | -876
farmers or forest workers | -876
rural areas | -876
myalgia | -168
fever | -168
thrombocytopenia | -168
month of August | -168
SFTS | 0
rhabdomyolysis | 0
acute febrile diseases | 0
leptospirosis | 0
human granulocytic anaplasmosis | 0
scrub typhus | 0
hemorrhagic fever renal syndrome | 0
co-infection | 0
seizure | -96
meningitis | -96
encephalitis | -96
spontaneous intracranial hemorrhage | -96
thrombocytopenia | -96
encephalitis or hemorrhage | 0
lumbar puncture | 0
electroencephalography | 0
prone position | 48
rapidly progressive acute respiratory distress syndrome | 48
multiple organ failure | 72
SFTS virus | 72
reverse transcriptase polymerase chain reaction | 72
Korea Centers for Disease Control and Prevention | 72
SFTS case reported in Korea | -876
SFTS cases reported | -876
farmers or forest workers | -876
rural areas | -876
myalgia | -168
fever | -168
thrombocytopenia | -168
month of August | -168
SFTS | 0
rhabdomyolysis | 0
acute febrile diseases | 0
leptospirosis | 0
human granulocytic anaplasmosis | 0
scrub typhus | 0
hemorrhagic fever renal syndrome | 0
co-infection | 0
seizure | -96
meningitis | -96
encephalitis | -96
spontaneous intracranial hemorrhage | -96
thrombocytopenia | -96
encephalitis or hemorrhage | 0
lumbar puncture | 0
electroencephalography | 0
prone position | 48
rapidly progressive acute respiratory distress syndrome | 48
multiple organ failure | 72
SFTS virus | 72
reverse transcriptase polymerase chain reaction | 72
Korea Centers for Disease Control and Prevention | 72
SFTS case reported in Korea | -876
SFTS cases reported | -876
farmers or forest workers | -876
rural areas | -876
myalgia | -168
fever | -168
thrombocytopenia | -168
month of August | -168
SFTS | 0
rhabdomyolysis | 0
acute febrile diseases | 0
leptospirosis | 0
human granulocytic anaplasmosis | 0
scrub typhus | 0
hemorrhagic fever renal syndrome | 0
co-infection | 0
seizure | -96
meningitis | -96
encephalitis | -96
spontaneous intracranial hemorrhage | -96
thrombocytopenia | -96
encephalitis or hemorrhage | 0
lumbar puncture | 0
electroencephalography | 0
prone position | 48
rapidly progressive acute respiratory distress syndrome | 48
multiple organ failure | 72
SFTS virus | 72
reverse transcriptase polymerase chain reaction | 72
Korea Centers for Disease Control and Prevention | 72
SFTS case reported in Korea | -876
SFTS cases reported | -876
farmers or forest workers | -876
rural areas | -876
myalgia | -168
fever | -168
thrombocytopenia | -168
month of August | -168
SFTS | 0
rhabdomyolysis | 0
acute febrile diseases | 0
leptospirosis | 0
human granulocytic anaplasmosis | 0
scrub typhus | 0
hemorrhagic fever renal syndrome | 0
co-infection | 0
seizure | -96
meningitis | -96
encephalitis | -96
spontaneous intracranial hemorrhage | -96
thrombocytopenia | -96
encephalitis or hemorrhage | 0
lumbar puncture | 0
electroencephalography | 0
prone position | 48
rapidly progressive acute respiratory distress syndrome | 48
multiple organ failure | 72
SFTS virus | 72
reverse transcriptase polymerase chain reaction | 72
Korea Centers for Disease Control and Prevention | 72
SFTS case reported in Korea | -876
SFTS cases reported | -876
farmers or forest workers | -876
rural areas | -876
myalgia | -168
fever | -168
thrombocytopenia | -168
month of August | -168
SFTS | 0
rhabdomyolysis | 0
acute febrile diseases | 0
leptospirosis | 0
human granulocytic anaplasmosis | 0
scrub typhus | 0
hemorrhagic fever renal syndrome | 0
co-infection | 0
seizure | -96
meningitis | -96
encephalitis | -96
spontaneous intracranial hemorrhage | -96
thrombocytopenia | -96
encephalitis or hemorrhage | 0
lumbar puncture | 0
electroencephalography | 0
prone position | 48
rapidly progressive acute respiratory distress syndrome | 48
multiple organ failure | 72
SFTS virus | 72
reverse transcriptase polymerase chain reaction | 72
Korea Centers for Disease Control and Prevention | 72
SFTS case reported in Korea | -876
SFTS cases reported | -876
farmers or forest workers | -876
rural areas | -876
myalgia | -168
fever | -168
thrombocytopenia | -168
month of August | -168
SFTS | 0
rhabdomyolysis | 0
acute febrile diseases | 0
leptospirosis | 0
human granulocytic anaplasmosis | 0
scrub typhus | 0
hemorrhagic fever renal syndrome | 0
co-infection | 0
seizure | -96
meningitis | -96
encephalitis | -96
spontaneous intracranial hemorrhage | -96
thrombocytopenia | -96
encephalitis or hemorrhage | 0
lumbar puncture | 0
electroencephalography | 0
prone position | 48
rapidly progressive acute respiratory distress syndrome | 48
multiple organ failure | 72
SFTS virus | 72
reverse transcriptase polymerase chain reaction | 72
Korea Centers for Disease Control and Prevention | 72
SFTS case reported in Korea | -876
SFTS cases reported | -876
farmers or forest workers | -876
rural areas | -876
myalgia | -168
fever | -168
thrombocytopenia | -168
month of August | -168
SFTS | 0
rhabdomyolysis | 0
acute febrile diseases | 0
leptospirosis | 0
human granulocytic anaplasmosis | 0
scrub typhus | 0
hemorrhagic fever renal syndrome | 0
co-infection | 0
seizure | -96
meningitis | -96
encephalitis | -96
spontaneous intracranial hemorrhage | -96
thrombocytopenia | -96
encephalitis or hemorrhage | 0
lumbar puncture | 0
electroencephalography | 0
prone position | 48
rapidly progressive acute respiratory distress syndrome | 48
multiple organ failure | 72
SFTS virus | 72
reverse transcriptase polymerase chain reaction | 72
Korea Centers for Disease Control and Prevention | 72
SFTS case reported in Korea | -876
SFTS cases reported | -876
farmers or forest workers | -876
rural areas | -876
myalgia | -168
fever | -168
thrombocytopenia | -168
month of August | -168
SFTS | 0
rhabdomyolysis | 0
acute febrile diseases | 0
leptospirosis | 0
human granulocytic anaplasmosis | 0
scrub typhus | 0
hemorrhagic fever renal syndrome | 0
co-infection | 0
seizure | -96
meningitis | -96
encephalitis | -96
spontaneous intracranial hemorrhage | -96
thrombocytopenia | -96
encephalitis or hemorrhage | 0
lumbar puncture | 0
electroencephalography | 0
prone position | 48
rapidly progressive acute respiratory distress syndrome | 48
multiple organ failure | 72
SFTS virus | 72
reverse transcriptase polymerase chain reaction | 72
Korea Centers for Disease Control and Prevention | 72
SFTS case reported in Korea | -876
SFTS cases reported | -876
farmers or forest workers | -876
rural areas | -876
myalgia | -168
fever | -168
thrombocytopenia | -168
month of August | -168
SFTS | 0
rhabdomyolysis | 0
acute febrile diseases | 0
leptospirosis | 0
human granulocytic anaplasmosis | 0
scrub typhus | 0
hemorrhagic fever renal syndrome | 0
co-infection | 0
seizure | -96
meningitis | -96
encephalitis | -96
spontaneous intracranial hemorrhage | -96
thrombocytopenia | -96
encephalitis or hemorrhage | 0
lumbar puncture | 0
electroencephalography | 0
prone position | 48
rapidly progressive acute respiratory distress syndrome | 48
multiple organ failure | 72
SFTS virus | 72
reverse transcriptase polymerase chain reaction | 72
Korea Centers for Disease Control and Prevention | 72
SFTS case reported in Korea | -876
SFTS cases reported | -876
farmers or forest workers | -876
rural areas | -876
myalgia | -168
fever | -168
thrombocytopenia | -168
month of August | -168
SFTS | 0
rhabdomyolysis | 0
acute febrile diseases | 0
leptospirosis | 0
human granulocytic anaplasmosis | 0
scrub typhus | 0
hemorrhagic fever renal syndrome | 0
co-infection | 0
seizure | -96
meningitis | -96
encephalitis | -96
spont