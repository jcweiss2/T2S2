45 years old | 0
African American | 0
male | 0
admitted to the hospital | 0
history of depression | -672
history of anxiety | -672
history of sleep disorder | -672
history of hypertension | -672
history of substance abuse | -672
elevated blood sugar | -336
methadone | -336
trazodone | -336
history of intravenous heroin abuse | -8760
history of inhalational cocaine abuse | -8760
abstinent from heroin and cocaine | -720
smoking cannabinoids | -13140
using K2 | -72
found unresponsive | 0
supply of K2 | 0
normal blood pressure | 0
tachycardia | 0
tachypnea | 0
high grade temperature | 0
hypoxia | 0
obtunded | 0
bilateral pupils equal and reactive to light | 0
normal tone | 0
absence of rigidity | 0
reflexes 1+ and symmetric | 0
no clonus | 0
no focal neurological deficits | 0
regular tachycardia | 0
marked hyperglycemia | 0
elevated creatinine | 0
hypernatremia | 0
hypokalemia | 0
severe hypophosphatemia | 0
mildly elevated cardiac enzymes | 0
hepatitis C Ab reactive | 0
HIV Ag/Ab non-reactive | 0
Ab reactivity to hepatitis A and hepatitis B Surface Ag | 0
sinus tachycardia | 0
first-degree atrioventricular block | 0
anion gap metabolic acidosis | 0
respiratory acidosis | 0
metabolic alkalosis | 0
hypertriglyceridemia | 0
subarachnoid hemorrhage | 0
possible parenchymal hemorrhage | 0
focal Fluid-attenuated inversion recovery (FLAIR) hyper-intense signal | 0
seizure prophylaxis | 24
improved mental status | 504
discharged | 504
STEMI | 24
reversible cardiomyopathy | 24
rhabdomyolysis | 24
severe metabolic derangement | 24
intubation for ventilator support | 24
hyperthermia | 0
no leukocytosis | 0
no bandemia | 0
afebrile | 24
negative blood and sputum culture | 48
negative urine analysis | 48
normal abdominal CT scan | 48
normal abdominal ultrasound | 48
new perihilar and bibasilar opacities | 72
broad-spectrum antibiotic therapy | 72
ampicillin sulbactam | 72
SIRS | 0
pneumonia | 72
normotensive | 0
elevated CPK | 0
peak CPK | 336
decreased CPK | 504
normal renal function | 504
positive urine toxicology for methadone | 0
negative toxicology screen for cannabinoids | 0
negative toxicology screen for flunitrazepam | 0
negative toxicology screen for gamma hydroxybutarate | 0
recovered entirely | 504