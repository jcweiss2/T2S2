73 years old | 0
female | 0
vaginal vault cancer stage 4 | -672
palliative RT to the vagina | -672
10 fractions of palliative RT | -672
1 cycle of chemotherapy | -672
shortness of breath | -168
fever | -168
constipation | -168
generalized weakness | -168
unresponsiveness | -168
admitted to the hospital | 0
oxygen saturation 89% on room air | 0
temperature 101.9F | 0
respiratory rate of 24 | 0
heart rate of 140 | 0
blood pressure measuring 110/65 | 0
purple urinary bag | -72
percutaneous nephrostomy (PCN) stents | -672
bilateral hydroureteronephrosis | -672
chronic kidney disease | -672
impingement of vaginal vault mass on both the ureters | -672
acute renal failure | -672
post-renal acute kidney failure | -672
Karnofsky performance status 40 | 0
colour change | -72
provisional diagnosis of PUBS | 0
high white blood cell count | 0
urinary pH 7.5 | 0
moderate leukocytes in the urine | 0
nitrates positive | 0
leucocyte esterase positive | 0
no ingestion of medications/food items | 0
no poisonous materials | 0
no haematuria | 0
no porphyria | 0
started on empirical IV cefoperazone and sulbactam | 0
started on levofloxacin 500 mg | 0
urine culture grew Escherichia coli | 0
urine culture grew Klebsiella spp. | 0
Gram-negative bacteremia | 0
urine discolouration subsided | 120
no clinical improvement | 120
disease burden | 120
ongoing sepsis | 120
multi-organ failure | 120
delirious | 144
increased breathlessness | 144
fever spikes | 144
condition deteriorated | 144
expired | 168