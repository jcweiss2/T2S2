52 years old | 0
male | 0
admitted to the hospital | 0
sore throat | -240
right laterocervical swelling | -240
diabetes | 0
no pharmacological allergies | 0
no psychosocial problems | 0
no family genetic disease | 0
inflammatory right laterocervical swelling | 0
trismus | 0
raised tongue | 0
right peritonsillar swelling | 0
bad dentition | 0
early signs of sepsis | 0
low-grade temperature | 0
mild tachycardia | 0
hemoglobin 13.2 g/dl | 0
WBC 13120/mm3 | 0
Absolute neutrophils 22530/mm3 | 0
C-reactive protein 441.9 mg/l | 0
creatinine 76.5 mg/L | 0
urea 0.69 g/L | 0
ASAT 585 UI/l | 0
ALAT 607 UI/l | 0
PT 48% | 0
fasting blood glucose 3.05 g/L | 0
multidrug-resistant streptococcus intermedius | 0
resistant to betalactamine | 0
resistant to tetracyclin | 0
resistant to ciprofloxacin | 0
resistant to erythromycin | 0
resistant to lincomycin | 0
resistant to trimethoprim/Sulfamethoxasol | 0
sensitive to levofloxacin | 0
sensitive to moxifloxacin | 0
sensitive to vancomycin | 0
thrombosed right IJV | 0
right tonsil abscess | 0
abscessed bilateral submandibular lymph nodes | 0
narrowing of the adjacent pharyngeal lumen | 0
emphisematous cervical cellulitis | 0
hospitalized | 0
multidisciplinary management | 0
broad-spectrum antibiotic therapy | -24
amoxicillin/clavulanic acid | 0
metronidazole | 0
gentamycin | 0
moxifloxacin | 96
anticoagulant therapy | 0
Enoxaparin | 0
Acenocoumarol | 96
endobucal adenophlegmon incision | 24
daily puncture of the right tonsil abscess | 0
increase in lateral cervical tumefaction | 48
emphysematous cervical facial cellulitis | 48
drainage of the collections | 72
sebileau incision | 72
cervical facial collections | 72
necrosis of the submandibular gland | 72
delbet drain | 72
communications closed | 72
good tolerance to the surgery | 96
good tolerance to post-operative care | 96
antibiotics | 0
local care | 0
no complications | 120
anticoagulated with heparin | 120
echocardiogram | 120
negative for endocarditis | 120
discharged | 288