64 years old | 0
male | 0
admitted to the hospital | 0
general malaise | 0
fever | 0
chills | 0
nuchal swelling | 0
facial swelling | 0
left-sided microtia | -259200
absence of meatus acusticus | -259200
diabetes mellitus type 2 | -6720
arterial hypertension | -6720
valsartan | -6720
head-and-neck edema | 0
herpetiform-grouped vesicles | 0
yellowish crusts | 0
bullae | 0
leukocytosis | 0
thrombocytopenia | 0
lowered hematocrit | 0
hemoglobin | 0
erythrocyte count | 0
neutrophilia | 0
lymphopenia | 0
increased number of large unstained cells | 0
C-reactive protein | 0
HIV tests | 0
antibiotic treatment with sultamicillin | 0
facial swelling worsened | 24
referred to Ear Nose Throat-department | 24
diagnostic ultrasound | 24
thoracic computerized tomography | 24
impetiginized herpes zoster | 48
antibiotic treatment changed to clindamycin | 48
aciclovir | 48
pain management with metamizole sodium | 48
minor clinical improvement | 72
blasts in peripheral blood | 72
bone marrow biopsy suggested | 72
bone marrow biopsy refused | 72
malodorous oozing | 96
formation of bullae | 96
increasing edema | 96
firm infiltrates | 96
skin biopsies | 96
histopathology | 96
putrid inflammation | 96
vesicles showed dissemination | 96
zoster generalisatus | 96
increased dosage of aciclovir | 120
pain sensations worsened | 120
pregabalin started | 120
certoparin sodium | 120
thrombosis prophylaxis | 120
CRP increased | 144
leukocytosis | 144
procalcitonin increased | 144
septicemia suspected | 144
transferred to intensive care unit | 144
central venous access | 144
subclavian catheter | 144
piperacillin | 144
levofloxacin | 144
acyclovir | 144
prednisolone | 144
doughy stool | 168
antibiosis changed to vancomycin | 168
stool samples for Clostridium difficile | 168
clinical improvement | 192
reduction of vesiculation | 192
reduction of edema | 192
CT | 192
bone marrow biopsy | 192
atypical myelopoiesis | 192
reduced atypical erythropoiesis | 192
micromegakaryocytic megakaryopoiesis | 192
bone marrow blasts | 192
myelodysplastic syndrome | 192
RAEB II | 192
chromosomal analysis | 192
cytodiagnostics | 192
karyotype 46/XY | 192
translocations t(2;12)(p13;q13) | 192
translocations t(6;9)(p22;q34) | 192
erythrocyte concentrates | 192
pain in right arm | 336
erythematous skin surrounding subclavian catheter | 336
catheter removed | 336
microbial cultures of catheter tip | 336
venous duplex sonography | 336
vena subclavia thrombosis | 336
soft tissue hematoma | 336
oozing of scalp | 360
oozing of ear helix | 360
microbial swaps | 360
Pseudomonas aeruginosa | 360
intensified diuresis | 360
progressive edema | 360
cytoreductive treatment with azacitidine | 360
anemia | 360
thrombocytopenia | 360
erythrocyte concentrates | 360
thrombocyte concentrates | 360
herpes zoster persisted | 360
varicella immunoglobulin | 384
anaphylactic shock | 384
septic shock | 408
death | 408