46 years old | 0
Asian-Indian | 0
male | 0
admitted to the hospital | 0
tropical chronic pancreatitis | -8760
oral pancreatic enzyme therapy | -8760
exocrine pancreatic insufficiency | -8760
non-insulin-dependent diabetes mellitus | -4380
glipizide | -4380
midepigastric pain | -6
epigastric pain | -6
pain control with narcotics | -6
discharged | -48
epigastric pain | -48
nausea | -48
vomiting | -48
CT scan | -48
fatty atrophy of pancreatic head | -48
fatty atrophy of uncinate process | -48
pancreatic duct filled with calcifications | -48
obstruction at the level of the neck | -48
upstream ductal dilatation | -48
admitted for management of pain | -48
chronic atrophic calcific pancreatitis | -144
dilated pancreatic duct | -144
intraductal calculi | -144
ERCP | -144
pancreatography | -144
medically managed | -144
discharged | -144
fever | 48
chills | 48
rigors | 48
severe sepsis | 48
septic shock | 48
transferred to intensive care unit | 48
intubated | 48
hypoxemic respiratory failure | 48
acute respiratory distress syndrome | 48
multiorgan failure | 48
broad-spectrum antibiotics | 48
vasopressor support | 48
activated recombinant human protein C | 48
ultrasound of abdomen | 48
dilated pancreatic duct | 48
calculus within the duct | 48
diffusely echogenic pancreas | 48
prominent common bile duct | 48
bedside emergency ERCP | 72
frank pus expelling through major papilla of Vater | 72
evacuation of pus | 72
cholangiogram | 72
pancreatogram | 72
guide wire introduced into pancreatic duct | 72
pus evacuated | 72
5-cm-long 5 F stent placed | 72
stent failed to show pus draining | 72
stent pulled out | 72
ASPD | 72
contrast enhanced CT scan | 96
inflammatory changes within fat surrounding pancreas | 96
edema | 96
diminished dilatation of pancreatic duct | 96
distal migration of calculus | 96
bilateral moderate pleural effusions | 96
clinical improvement | 96
stabilization of hemodynamic parameters | 96
blood cultures grew Klebsiella ornithinolytica | 96
extubated | 120
transferred from intensive care unit | 120
completed antibiotic course | 120
discharged home | 264
follow-up examinations | 720
follow-up examinations | 2160
no further complications | 720
no further complications | 2160