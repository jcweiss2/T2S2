Here is the table of events and timestamps:

57 years old | 0
Hispanic | 0
history of coronary artery disease | -2160
myocardial infarction | -2160
ischemic dilated cardiomyopathy | -2160
pocket infection of his cardiac resynchronization therapy defibrillator | -144
cardiac resynchronization therapy defibrillator | -2160
generator change | -144
erythema and discomfort around his left upper chest implant site | -672
edema and serosanguinous drainage | -672
oral amoxicillin treatment | -672
nonbacteremic | -144
afebrile | -144
laboratory investigations within normal limits | -144
echocardiography severely reduced left ventricular systolic function | -144
ejection fraction 20%–25% | -144
global hypokinesis of the left ventricle | -144
no evidence of vegetations | -144
preoperative computed tomography leads scarred to the lateral wall of the superior vena cava | -144
transvenous lead extraction | 0
device removed | 0
coronary sinus and right atrial leads extracted | 0
hypotensive | -1
transesophageal echocardiography large pericardial effusion | -1
emergency midsternotomy | -1
5-mm tear in the superior cavoatrial junction | -1
perforation in the right atrium | -1
oozing hematoma at the level of the innominate vein | -1
bleeding manually controlled with pressure | -1
cardiopulmonary bypass instituted | -1
right ventricular lead capped and abandoned | -1
intra-aortic balloon pump placed | -1
multiple blood transfusions | -1
coagulopathy | -1
cryoprecipitate transfusions | -1
platelets transfusions | -1
fresh frozen plasma transfusions | -1
factor VII transfusions | -1
chest closed | -1
26 units of blood products given intraoperatively | -1
10 units of packed red blood cells given intraoperatively | -1
postoperative transfer to the intensive care unit | -1
severe cardiogenic shock | -1
multiorgan failure | -1
hypotensive | -1
large doses of vasopressin | -1
epinephrine | -1
norepinephrine | -1
hypoxic respiratory failure | -1
mechanical ventilation | -1
liver failure | -1
albumin given | -1
continuous venovenous hemodialysis | -1
bilateral, symmetrical cyanotic changes to all 5 digits of his upper and lower extremities | -1
vasopressor administration stopped | -1
upper- and lower-digit ischemia progressed to dry gangrene | -9
dull pain | -9
inability to move fingers and toes | -9
bilateral stiffness | -9
2+ pitting edema | -9
nonexistent capillary refill time | -9
palpable 2+ peripheral pulses | -9
Doppler study flat waveforms on all digits and toes bilaterally | -9
no proximal occlusion or stenosis | -9
intra-aortic balloon pump removed | 7
endotracheal tube removed | 7
albumin discontinued | 11
liver enzymes returned to normal limits | 11
kidney function gradually improved | 41
hemodialysis stopped | 41
mental status improved | 41
necrotic lesions treated conservatively | 41
povidone-iodine dressings | 41
debridement | 27
negative-pressure wound therapy | 27
purulent, foul-smelling material from his left infraclavicular operative site | 27
stabilized and transferred to our facility | 54
preoperative transesophageal echocardiography | 54
diminished ejection fraction 10%–15% | 54
laser extraction of his retained lead | 58
pus drained from the subfascial area | 58
appropriate antibiotic regimen | 58
transesophageal echocardiography | 58
implantable cardioverter-defibrillator system implanted | 64
evaluation of his hands and feet | 64
no signs of local infection or wet gangrene | 64
black skin changes and demarcation lines | 64
frank mummification of his digits and toes | 64
discharged to home health services | 77
amputation and debridement of his necrotic feet | 106
amputation of his fingers scheduled | 106