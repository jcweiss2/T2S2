54 years old | 0
    non-smoking | 0
    woman | 0
    stage IV lung adenocarcinoma | 0
    brain metastasis | 0
    liver metastasis | 0
    multiple bone metastasis | 0
    ECOG score 0 | 0
    chronic cough | 0
    CT-guided biopsy of right lung tumor | 0
    L858R-positive lung adenocarcinoma | 0
    clinical staging cT4N3M1b | 0
    disease progression | -175200
    erlotinib use | -175200
    osimertinib use | -157680
    chemotherapy | -126576
    disease progression | -7008
    re-biopsy at right middle lobe | -7008
    genomic profiling | -7008
    ACTDrug NGS-based assay | -7008
    mutations L858R/cis-T790M/cis-C797S | -7008
    no other molecular alterations | -7008
    brigatinib use | 0
    afatinib combination suggested | 0
    off-label treatment agreement | 0
    brigatinib 90 mg once daily | 0
    afatinib 30 mg once daily | 0
    admission | 0
    exertional dyspnea | 48
    dry cough | 48
    hypercapnic respiratory failure | 72
    intubation | 72
    leukocytosis | 72
    neutrophil predominant | 72
    carbon dioxide retention | 72
    bilateral interstitial infiltrates | 72
    pneumonia | 72
    broad-spectrum antibiotics | 72
    fever subsided | 72
    septic shock improvement | 72
    poor oxygenation | 72
    bilateral ground-glass opacities | 72
    left lower lung consolidation | 72
    negative microbiology studies | 72
    EOPEs of doubled tyrosine kinase inhibitors | 72
    intravenous methylprednisolone 40 mg every 8 hours | 72
    oxygenation improvement | 120
    bilateral infiltrates improvement | 120
    complete resolution of ground-glass opacities | 336
    complete resolution of consolidation | 336
    transfer to respiratory care center | 504
    weaning | 504
    intensive care unit transfer | 504
    seizure due to brain metastasis | 504
    brain radiotherapy | 504
    progressive septic shock | 504
    broad-spectrum antibiotics | 504
    vasopressors | 504
    death | 864
    
    