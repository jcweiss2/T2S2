34 years old | 0
    multipara | 0
    visited the ER | 0
    low abdominal pain | 0
    nausea | 0
    vomiting | 0
    157 cm in height | 0
    weighed 67 kg | 0
    weight gain during pregnancy | 0
    parity 1-0-0-1 | 0
    no abnormalities in past medical history | 0
    blood pressure 120/75 mmHg | 0
    heart rate 75 beats/min | 0
    respiratory rate 22 times/min | 0
    chest radiography normal | 0
    ST segment depression | 0
    troponin-T increased to 0.206 ng/ml | 0
    CK-MB 3.52 ng/ml | 0
    no other lab abnormalities | 0
    fetal heart rate 130 beats/min | 0
    blood pressure increased to 158/100 mmHg | 1
    sinus tachycardia 124 beats/min | 1
    left ventricle size normal | 1
    moderate decline in systolic function | 1
    decrease in overall wall motion | 1
    moderate mitral regurgitation | 1
    tricuspid regurgitation | 1
    pulmonary hypertension | 1
    LVEF 39% | 1
    LVEDD 5.2 cm | 1
    LVESD 4.3 cm | 1
    transferred to intensive care | 1
    blood pressure 149/100 mmHg | 1
    heart rate 110 beats/min | 1
    respiration rate 27 times/min | 1
    hemoptysis | 4
    dyspnea | 4
    oxygen via nasal prong 4 L/min | 4
    chest radiograph severe pulmonary edema | 4
    furosemide 20 mg | 4
    nitroglycerin 8 µg/min | 4
    no improvement | 4
    additional furosemide 20 mg | 4
    nitroglycerin increased to 12 µg/min | 4
    oxygen via mask 10 L/min | 4
    ABGA pH 7.4 | 4
    PaCO2 16.1 mmHg | 4
    PaO2 62 mmHg | 4
    BE -8.7 mEq/L | 4
    SaO2 91% | 4
    fetal heart rate 180 beats/min | 4
    fetal distress anticipated | 4
    cesarean section decided | 4
    severe dyspnea | 4
    orthopnea | 4
    hemoptysis worsened when lying down | 4
    blood pressure 130/98 mmHg | 4
    heart rate 128 beats/min | 4
    respiratory rate 45 times/min | 4
    sinus tachycardia | 4
    general anesthesia for cesarean section | 4
    ECMO attempted | 4
    ECMO installation failed | 4
    ECMO under general anesthesia | 4
    arrived at operating room | 4
    oxygen 10 L/min via mask | 4
    nitroglycerin 12 µg/min | 4
    ECG monitoring | 4
    noninvasive blood pressure monitor | 4
    pulse oximeter | 4
    catheter in right radial artery | 4
    blood pressure 135/98 mmHg | 4
    heart rate 130 beats/min | 4
    peripheral oxygen saturation 98% | 4
    ABGA pH 7.40 | 4
    PaCO2 22 mmHg | 4
    PaO2 82 mmHg | 4
    BE -9.3 mEq/L | 4
    SaO2 96% | 4
    blood pressure 140/105 mmHg | 4
    heart rate 132 beats/min | 4
    thiopental sodium 250 mg | 4
    succinylcholine 100 mg | 4
    intubation | 4
    atracurium 40 mg | 4
    sevoflurane 2 vol% | 4
    tidal volume 550 ml | 4
    respiration rate 16 times/min | 4
    PEEP 5 cmH2O | 4
    blood pressure 155/110 mmHg | 4
    heart rate 138 beats/min | 4
    sinus tachycardia | 4
    ABGA pH 7.39 | 4
    PaCO2 24 mmHg | 4
    PaO2 70 mmHg | 4
    BE -9.2 mEq/L | 4
    SaO2 93% | 4
    ECMO applied | 4
    femoral arterial cannula | 4
    femoral venous cannula | 4
    ECMO installation time 20 minutes | 4
    flow rate 3 L/min | 4
    central venous catheter inserted | 4
    Swan-Ganz catheter attempted | 4
    Swan-Ganz catheter advanced to right ventricle | 4
    blood pressure 140-160/100-110 mmHg | 4
    heart rate 120-130 beats/min | 4
    peripheral oxygen saturation 91-95% | 4
    central venous pressure 22-24 mmHg | 4
    tidal volume adjusted to 400 ml | 4
    respiration rate 10 times/min | 4
    FiO2 0.5 | 4
    nitroglycerin continued | 4
    infant delivered | 4
    APGAR scores 3 and 4 | 4
    infant intubation | 4
    oxytocin 40 units | 4
    colloid solution 500 ml | 4
    blood pressure mean 100-120 mmHg | 4
    heart rate 100 beats/min | 4
    peripheral oxygen saturation 100% | 4
    central venous pressure 14-18 mmHg | 4
    ABGA pH 7.38 | 4
    PaCO2 24.6 mmHg | 4
    PaO2 408 mmHg | 4
    BE -11 mEq/L | 4
    SaO2 100% | 4
    operating time 1 hour 40 minutes | 4
    anesthetic time 1 hour 45 minutes | 4
    blood loss 1000 ml | 4
    fluid volume 600 ml | 4
    transferred to ICU | 4
    ECMO maintained | 4
    intubation maintained | 4
    blood pressure 90-100 mmHg | 4
    heart rate 110 beats/min | 4
    peripheral oxygen saturation 100% | 4
    ABGA pH 7.31 | 4
    PaCO2 22 mmHg | 4
    PaO2 359 mmHg | 4
    BE -13.2 mEq/L | 4
    SaO2 100% | 4
    ECMO flow decreased to 2 L/min | 72
    blood pressure 95-120/79-95 mmHg | 72
    heart rate 90-110 beats/min | 72
    peripheral oxygen saturation 100% | 72
    central venous pressure 5-8 mmHg | 72
    ABGA pH 7.5 | 72
    PaCO2 28 mmHg | 72
    PaO2 508 mmHg | 72
    BE 0.8 mEq/L | 72
    SaO2 100% | 72
    tidal volume 400 ml | 72
    respiration rate 12 times/min | 72
    PEEP 3 cmH2O | 72
    FiO2 0.4 | 72
    ECMO flow decreased to 1.3 L/min | 96
    blood pressure 120-140/90-100 mmHg | 96
    heart rate 90-100 beats/min | 96
    peripheral oxygen saturation 100% | 96
    central venous pressure 4-8 mmHg | 96
    ABGA pH 7.48 | 96
    PaCO2 32 mmHg | 96
    PaO2 517 mmHg | 96
    BE 0.6 mEq/L | 96
    SaO2 100% | 96
    ECMO flow decreased to 1 L/min | 108
    blood pressure 110-140/80-100 mmHg | 120
    heart rate 80-100 beats/min | 120
    peripheral oxygen saturation 100% | 120
    central venous pressure 9 mmHg | 120
    ABGA pH 7.54 | 120
    PaCO2 28 mmHg | 120
    PaO2 639 mmHg | 120
    BE 1.8 mEq/L | 120
    SaO2 100% | 120
    ECMO removed | 120
    blood pressure 94-104/66-70 mmHg | 120
    heart rate 100 beats/min | 120
    peripheral oxygen saturation 100% | 120
    central venous pressure 5-7 mmHg | 120
    ABGA pH 7.4 | 120
    PaCO2 28 mmHg | 120
    PaO2 639 mmHg | 120
    BE 1.8 mEq/L | 120
    SaO2 100% | 120
    dopamine 5 µg/kg/min | 120
    mechanical ventilation removed | 168
    transferred to general ward | 168
    blood pressure 100-130/65-70 mmHg | 168
    heart rate 75-90 beats/min | 168
    ABGA pH 7.42 | 168
    PaCO2 43 mmHg | 168
    PaO2 156 mmHg | 168
    BE 2.9 mEq/L | 168
    SaO2 98% | 168
    ECG normal | 168
    pulmonary edema improved | 168
    LVEF 58% | 168
    slight mitral regurgitation | 168
    infant transferred to NICU | 4
    babygram normal | 24
    extubation after 2 days | 48
    abdominal sonography normal | 48
    brain MRI no ischemia | 48
    infant discharged after 11 days | 264