63 years old | 0
male | 0
admitted to the hospital | 0
productive cough | -48
dyspnea | -48
pulmonary tuberculosis | -8760
smoking | -8760
mediastinal enlargement | 0
bulging on the right atrium contour | 0
afebrile | 0
normal hemodynamic parameters | 0
no peripheral edema | 0
normal lung examination | 0
ejection murmur | 0
raised jugular venous pressure | 0
hepatomegaly | 0
pericardium thickening | 0
mild effusion | 0
left ventricular ejection fraction of 60% | 0
mass with soft tissue attenuation | 0
infiltrating the pericardium | 0
infiltrating the anterior wall of the right atrium | 0
multiple, bilateral, scattered, solid pulmonary nodules | 0
mass with heterogeneous distinction | 0
diffusely involving the pericardium | 0
compression/invasion of the right ventricle’s outflow tract | 0
compression/invasion of the pulmonary artery | 0
compression/invasion of the superior vena cava | 0
pericardium biopsied | 0
no evidence of malignancy | 0
pulmonary nodule biopsied | 0
mesenchymal malignancy | 0
sinusoidal vascular channels filled with red blood cells | 0
atypical endothelial cells | 0
positivity for CD31 | 0
positivity for CD34 | 0
negativity for Desmin | 0
negativity for S100 Protein | 0
diagnosis of angiosarcoma | 0
metastatic angiosarcoma | 0
primary to the right atrium | 0
chemotherapy with doxorubicin | 0
chemotherapy with ifosfamide | 0
reduction in the size of the pulmonary nodules | 504
pulmonary infection | 1008
refractory septic shock | 1032
death | 1056