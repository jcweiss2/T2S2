16 years old | 0
male | 0
admitted to the hospital | 0
severe fatigue | -672
computed tomography | -672
anterior mediastinal tumor | -672
hepatosplenomegaly | -672
lymph node swelling | -672
T-lymphoblastic lymphoma | -672
treated with cytotoxic agents | -672
Eastern Cooperative Oncology Group performance status 1 | 0
mild hepatosplenomegaly | 0
electrocardiogram normal | 0
serum brain natriuretic peptide 17.2 pg/mL | 0
transthoracic echocardiography normal | 0
left ventricular ejection fraction 59.8% | 0
induction treatment | -672
cyclophosphamide 750 mg/m2 | -672
doxorubicin 50 mg/m2 | -672
vincristine 2 mg/body | -672
prednisolone 60 mg/m2 | -672
L-asparaginase 6,000 U/m2 | -672
intrathecal injection | -672
consolidation treatment | -504
cyclophosphamide 750 mg/m2 | -504
therarubicin 25 mg/m2 | -504
cytarabine 75 mg/m2 | -504
6-mercaptoprine 50 mg/m2 | -504
intrathecal injection | -504
sanctuary treatment | -336
methotrexate 3,000 mg/m2 | -336
intrathecal injection | -336
re-induction treatment | -210
prednisolone 90 mg/m2 | -210
daunorubicin 50 mg/m2 | -210
cyclophosphamide 750 mg/m2 | -210
vincristine 2 mg/body | -210
L-asparaginase 5,000 U/body | -210
etoposide 100 mg/m2 | -210
bridging to conditioning | -126
doxorubicin 40 mg/m2 | -126
cyclophosphamide 500 mg/m2 | -126
vincristine 2 mg/body | -126
radiation 20 Gy/10 fr | -126
conditioning regimen | 0
etoposide 15 mg/kg | -10
cyclophosphamide 60 mg/kg | -8
total body irradiation 12 Gy/6 fr | -3
cord blood cell transplantation | 0
fever 38.6°C | -96
meropenem | -96
fever resolved | -92
high fever | 48
septic shock | 72
vancomycin | 72
transferred to intensive-care unit | 72
circulatory assisting agents | 72
respiratory condition worsened | 144
mechanical ventilation | 144
left ventricular ejection fraction 10.3% | 144
acute heart failure | 144
left ventricular wall thickness | 144
electrocardiogram abnormal | 144
R wave voltage 0.44 mV | 216
methylprednisolone 1.2 mg/kg/day | 216
body temperature 38-41°C | 216
dobutamine dose increased | 216
milrinone added | 216
cardiac exhaustion | 216
ivabradine 5 mg/day | 312
heart rate decreased | 312
dobutamine dose reduced | 312
BNP level decreased | 312
carvedilol 1.25 mg/day | 352
ivabradine dose increased | 352
carvedilol dose increased | 352
dobutamine and milrinone ceased | 424
discharged from ICU | 424
ventilator withdrawn | 504
engraftment recognized | 228
neutrophils | 228
red blood cells | 336
platelets | 384
grade 3 acute graft-versus-host disease | 336
methylprednisolone 2 mg/kg/day | 336
serum troponin I concentration decreased | 336
LVEF improved | 648
ECG improved | 648
R wave voltage 1.53 mV | 648
died of relapsed lymphoma | 1008