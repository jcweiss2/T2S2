59 years old | 0
female | 0
admitted to the hospital | 0
fever | -120
cough | -120
nasal obstruction | -120
diarrhea | -120
hypertension | -120
diabetes | -120
axillary temperature 38.5°C | 0
blood pressure 170/102 mm Hg | 0
respiratory rate 20 breaths per minute | 0
oxygen saturation 93% | 0
leukocytes 9260 per microliter | 0
D-dimer 2404 ng/mL | 0
fibrinogen 954 mg/dL | 0
SARS-CoV-2 positive | 0
ground-glass opacities in both lungs | 0
ceftriaxone | 0
azithromycin | 0
oseltamivir | 0
prophylactic low molecular weight heparin | 0
supplemental oxygen | 0
tachypnea | 24
dyspnea at rest | 24
oxygen saturation decreased to 88% | 24
intubation | 24
mechanical ventilation | 24
fibrinogen 729 mg/dL | 24
interleukin (IL)-6 149 | 24
antithrombin III 107% | 24
D-dimer 40,130 ng/mL | 24
pulmonary thromboembolism | 24
low molecular weight heparin 1 mg/kg twice daily | 24
CT angiography of the chest | 24
signs of acute pulmonary thromboembolism | 24
extubation | 168
pain in the right lower limb | 192
right second toe turned blue | 192
acute arterial occlusion | 192
femoral arterial line removal | 192
venous Doppler of the lower limbs | 192
transthoracic echocardiogram | 192
mild tricuspid regurgitation | 192
Right Ventricular Systolic Pressure of 40 mm Hg | 192
arteriography | 192
significant stenosis in posterior tibial artery | 192
tibiofibular trunk | 192
fibular artery | 192
angioplasty of the right lower limb | 192
amputation of the right second toe | 216
discharged from the hospital | 216
Apixaban 5 mg twice a day | 216
follow-up at the vascular surgeon’s office | 360
amputation stump in great condition | 360
no new complaints | 360
no respiratory symptoms | 360