82 years old| 0
female | 0
admitted to the emergency department | 0
hematemesis | 0
upper gastrointestinal bleeding suspicion | 0
decreased hemoglobin | 0
elevated infection signs | 0
leukocyte count 27 × 10^9/L | 0
C-reactive protein 15 mg/dL |; 0
soft abdomen | 0
diffuse tenderness | 0
no voluntary guarding | 0
beginning septic shock | 0
increasing hemodynamic instability | 0
loss of vigilance | 0
referred to intensive care unit | 0
intubation | 0
gastroscopy | 0
no upper gastrointestinal bleeding | 0
gallbladder penetration | 0
gallstones in the duodenal bulb | 0
computed tomography confirmation | 0
chronic cholecystitis | 0
pneumobilia | 0
gallbladder penetration in the duodenal bulb | 0
entry of gallstones in the intestine | 0
reflective intestinal atony | 0
dilated stomach | 0
filled with contrast medium | 0
Bouveret syndrome diagnosis | 0
sepsis | 0
open cholecystectomy | 0
gallstone salvage from the duodenum | 0
no biliary enteric fistula | 0
diabetes | 0
arterial hypertension | 0
no history of biliary symptoms | 0
discharged | 120
