60 years old | 0
male | 0
biopsy proven PAN | -8760
paroxysmal atrial fibrillation | -8760
hypertension | -8760
dyslipidemia | -8760
non-insulin dependent diabetes mellitus | -8760
admission for septic shock | -8760
scrotal pain | 0
fever | 0
103°F | 0
tachycardic | 0
130 beats per minute | 0
hypotensive | 0
103/40 mm Hg | 0
broad-spectrum antibiotics | 0
vancomycin | 0
Zosyn | 0
admission under medicine service | 0
kidney function worsened | 24
switch in antibiotics | 24
meropenem | 24
creatinine level continued to rise | 48
macular rash | 168
axillary area | 168
chest | 168
head | 168
neck | 168
abdomen | 168
decline of mental status | 168
worsening of skin lesions | 168
bullae | 168
vesicles | 168
dermatology team | 168
biopsy | 168
local steroid cream | 168
AGEP | 168
kidney injury | 168
neutrophilia | 168
cyclic fevers | 168
rash became pustular | 216
high grade fever | 216
109°F | 216
transfer to the intensive care unit | 216
cooling | 216
pulse steroids | 216
fever subsided | 240
improvement of the initial rash | 240
decreased progression of sloughing | 240
complete resolution of acute kidney injury | 240
taper in steroids | 240
intra- and subcorneal spongiform | 0
superficial, interstitial, mid-dermal infiltrate rich in neutrophils | 0
dermal edema | 0
discharged | 336