65 years old | 0
female | 0
admitted to the hospital | 0
recurrent fever | -720
nausea | -168
vomiting | -168
highest body temperature 38 ℃ | -720
neutrophil count 6.96×10^9/L ↑ | 0
monocyte count 0.86×10^9/L ↑ | 0
lymphocyte percentage 14.9% ↓ | 0
red blood cell count 3.17×10^12/L ↓ | 0
hemoglobin content 87 g/L ↓ | 0
hematocrit 0.28 L/L ↓ | 0
average red blood cell hemoglobin concentration 312 g/L ↓ | 0
platelet count 363×10^9/L ↑ | 0
platelet distribution width 8.3 fl ↓ | 0
C-reactive protein (CRP) 52.01 mg/L ↑ | 0
diagnosed with secondary infectious thrombocytopenia | 0
diagnosed with gram-negative bacilli septicemia (Klebsiella pneumoniae) | 0
diagnosed with liver abscess | 0
diagnosed with bilateral lung inflammation | 0
diagnosed with type 2 diabetes | 0
diagnosed with hypertension grade 3 (extremely high risk) | 0
given vancomycin | 0
given caspofungin | 0
given dexamethasone | 0
given posaconazole oral suspension | 0
liver abscess puncture and drainage treatment | 24
inflammatory indexes decreased | 48
light perception disappeared in the left eye | 72
eyelid redness and pain | 72
purulent secretion | 72
repeated fever | 72
left-sided headache | 72
diagnosed with endogenous endophthalmitis (left) | 72
diagnosed with orbital cellulitis (left) | 72
diagnosed with rubeosis iridis (left) | 72
diagnosed with exudative retinal detachment (left) | 72
diagnosed with diabetic retinopathy (right) | 72
intravitreal injection with vancomycin and ceftazidime | 72
symptoms relieved | 96
systemic infection under control | 96
left eyeball enucleation | 168
fever again after the operation | 168
given moxifloxacin | 168
given sulperazon | 168
temperature elevated again | 192
CT examination | 192
inflammation of both lungs | 192
pericardial effusion | 192
bilateral pleural thickening and effusion | 192
atelectasis in right inferior lobe | 192
liver cyst | 192
liver abscess | 192
right renal cyst | 192
myoma of the uterus | 192
history of hypertension | -8760
highest blood pressure 180/100 mmHg | -8760
oral valsartan | -8760
blood pressure controlled at 140/80 mmHg | -8760
no special history of other systematic diseases | 0
no history of surgery | 0
no history of blood transfusion | 0
no history of drug allergy | 0
diagnosed with sepsis | 0
diagnosed with secondary thrombocytopenia | 0
diagnosed with liver abscess | 0
diagnosed with gram-negative bacilli sepsis (Klebsiella pneumoniae) | 0
diagnosed with infection of lumbar vertebrae | 0
diagnosed with mesenteric panniculitis | 0
diagnosed with pelvic effusion | 0
diagnosed with pericardial effusion | 0
diagnosed with suppurative endophthalmitis (left) | 0
diagnosed with orbital cellulitis (left) | 0
diagnosed with retinal detachment (left) | 0
diagnosed with choroidal detachment (left) | 0
diagnosed with type 2 diabetes retinopathy (right) | 0
diagnosed with cortical senile cataract (right, immature stage) | 0
diagnosed with type 2 diabetes | 0
diagnosed with type 2 diabetes nephropathy stage I | 0
diagnosed with type 2 diabetic peripheral neuropathy | 0
diagnosed with hypertension grade 3 (extremely high risk) | 0
diagnosed with hepatic cyst | 0
diagnosed with renal cyst | 0
diagnosed with hypoproteinemia | 0
diagnosed with coronary atherosclerotic heart disease | 0
diagnosed with lacunar cerebral infarction | 0
diagnosed with moderate anemia | 0
diagnosed with risk of malnutrition | 0
convulsion with unconsciousness | 240
transferred to the respiratory intensive care unit | 240
CT examination | 240
lacunar infarction | 240
encephalomalacia | 240
bilateral pleural effusion | 240
lower lobe of the right lung insufficiently inflated | 240
intracranial infection | 240
lumbar puncture | 240
cerebrospinal fluid (CSF) analysis | 240
microbial metagenomic next-generation sequencing (mNGS) | 240
biochemistry analysis | 240
glucose <1.1 mmol/L ↓ | 240
chlorine 108 mmol/L ↓ | 240
CSF protein >3,000 mg/L ↑ | 240
mNGS results showed high sequence of Klebsiella pneumoniae with drug-resistant gene blaSHV | 240
given 2 g meropenem q8h prolonged for 3 hours | 240
body temperature improved | 264
blood routine improved | 264
CRP improved | 264
CT examination | 336
pulmonary edema and pleural effusion dissipated and absorbed | 336
CSF analysis | 336
chlorine 119 mmol/L ↓ | 336
micro amount of proteins 1,107 mg/L ↑ | 336
microalbumin 816.3 mg/L ↑ | 336
immunoglobulin G 308.5 mg/L ↑ | 336
α2-macroglobulin 18.5 mg/L ↑ | 336
β2-microglobulin 2.67 mg/L ↑ | 336
discharged from the hospital | 432