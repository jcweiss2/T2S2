67 years old | 0 | 0 
female | 0 | 0 
admitted to the hospital | 0 | 0 
backache | -24 | 0 
calculi in both kidneys | -24 | 0 
ureteral calculi | -24 | 0 
HLL | -0.5 | 0 
double J catheterization | -0.5 | 0 
purulent urine | -0.5 | 0 
fever | 0 | 48 
chill | 0 | 48 
low blood pressure | 0 | 48 
imipenem and Cilastatin sodium | 0 | 48 
fluid resuscitation | 0 | 48 
Norepinephrine | 0 | 48 
Hydrocortisone sodium succinate | 0 | 48 
anuria | 48 | 120 
ARDS | 48 | 120 
invasive ventilatory support | 48 | 120 
CRRT | 48 | 120 
transfer to ICU | 48 | 48 
sedated state | 48 | 48 
blood pressure 80/62 mmHg | 48 | 48 
heart rate 139 beats/min | 48 | 48 
transcutaneous oxygen saturation 80% | 48 | 48 
cold, clammy extremities | 48 | 48 
loud bubbling sound in the lung | 48 | 48 
arterial blood gas analysis | 48 | 48 
lactic acid 10.6 mmol/L | 48 | 48 
bicarbonate 10.8 mmol/L | 48 | 48 
central venous pressure 20 cmH2O | 48 | 48 
B lines in lung ultrasonography | 48 | 48 
diffuse dysfunction in left ventricle | 48 | 48 
LVEF 20.3% | 48 | 48 
sinus tachycardia | 48 | 48 
broad ST depression | 48 | 48 
elevated troponin I | 48 | 48 
elevated amino-terminal brain natriuretic peptide precursor | 48 | 48 
creatinine 356 μmol/L | 48 | 48 
VA-ECMO | 48 | 144 
CRRT | 48 | 144 
imipenem and Cilastatin sodium and Vancomycin | 48 | 120 
Norepinephrine stopped | 78 | 78 
Epinephrine stopped | 78 | 78 
lactic acid level declined | 90 | 90 
vasoactive drugs stopped | 138 | 138 
arterial blood lactate level normal | 144 | 144 
extended-spectrum β-lactamase-positive Escherichia coli | 48 | 48 
inflammatory indices diminished | 120 | 120 
anti-infection regimen continued | 120 | 240 
minimum serum trough concentration of Vancomycin monitored | 120 | 240 
LVEF 35% | 120 | 120 
necrotic skin | 120 | 120 
ECMO therapy weaned | 144 | 144 
CRRT discontinued | 144 | 144 
renal function scaled as acute kidney injury grade 3 | 144 | 144 
urine volume increased | 144 | 240 
vascular ultrasonography and computed tomography angiography | 240 | 240 
vascular surgery consultation | 240 | 240 
necrotic tissues amputated | 336 | 336 
tracheal intubation | 48 | 240 
spontaneous breathing | 120 | 120 
tracheotomy | 240 | 240 
anti-infective therapy replaced | 240 | 240 
physical rehabilitation | 240 | 240 
ventilator weaned | 480 | 480 
tracheotomy tube sealed | 600 | 600 
discharged | 768 | 768 
intermittent hemodialysis | 768 | 888 
self-care | 888 | 888 
intermittent hemodialysis continued | 888 | 888