38 years old | 0
female | 0
abdominal pain | 0
polyuria | 0
polydipsia | 0
nausea | 0
vomiting | 0
blood pressure 93/53 mmHg | 0
pulse 119 beats/min | 0
respiratory rate 28 breaths/min | 0
oxygen saturation 99% | 0
temperature 97.8°F | 0
Kussmaul breathing | 0
normal cardiopulmonary auscultation | 0
soft abdomen | 0
non-tender abdomen | 0
alert | 0
oriented | 0
blood pH 6.98 | 0
serum bicarbonate 5mmol/L | 0
serum anion gap 22 | 0
normal serum lactate | 0
serum glucose 506mg/dL | 0
urinalysis positive for ketones | 0
urine pregnancy test negative | 0
portable chest radiograph interstitial prominence | 0
portable chest radiograph ill-defined nodular opacities | 0
intravenous crystalloid 4 liters | 0
insulin infusion | 0
blood cultures collected | 0
admitted to intensive care unit | 0
hypoxemic | 0
dyspneic | 0
non-rebreather mask | 0
temperature 104°F | 0
obtundation | 0
diffuse crackles | 0
endotracheal intubation | 0
hypoxemic respiratory failure | 0
volume assist-control ventilation | 0
repeat chest radiograph diffuse bilateral opacities | 0
PaO2 59 mmHg | 0
PaO2/FiO2 ratio 84 | 0
lung-protective ventilation | 0
tidal volume 350ml | 0
PEEP 7.5 cmH2O | 0
vancomycin | 0
piperacillin/tazobactam | 0
blood cultures gram negative bacilli | 0
imipenem | 0
hemodynamic deterioration | 0
high-dose norepinephrine infusion | 0
vasopressin | 0
FiO2 100% | 24
PEEP 15 cmH2O | 24
inhaled nitric oxide therapy | 24
Klebsiella pneumoniae identification | 24
ceftriaxone | 24
abdominal ultrasonography | 24
complex avascular hepatic mass-like lesion | 24
interventional radiology drainage catheter | 24
pulseless electrical activity | 24
cardiopulmonary resuscitation | 24
resuscitative efforts aborted | 24
patient expired | 24
autopsy liver abscess | 24
lung sections diffuse abscess formation | 24
hyaline membranes | 24
diffuse alveolar damage | 24
invasive KLA syndrome | 24
ARDS | 24
