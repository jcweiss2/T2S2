72 years old | 0
male | 0
admitted to the hospital | 0
fever | -168
non-productive cough | -168
shortness of breath | -168
positive SARS-CoV-2 PCR test | -168
respiratory rate 55 breaths per minute | 0
peripheral oxygen saturation 74% | 0
oxygen therapy with non-rebreather mask | 0
blood pressure 144/91 mmHg | 0
heart rate 145 beats per minute | 0
body temperature 36.8°C | 0
increased white cell count | 0
lymphocytes 8% | 0
normal platelet count | 0
blood gas analysis | 0
pH 7.42 | 0
pCO2 23 mmHg | 0
pO2 43 mmHg | 0
HCO3 15 mmol/L | 0
base deficit -9 mmol/L | 0
lactic acid 7.46 mmol/L | 0
blood urea nitrogen 36 mg/dL | 0
creatinine 1.4 mg/dL | 0
alanine aminotransferase 169 U/L | 0
aspartate aminotransferase 238 U/L | 0
procalcitonin 51.36 ng/mL | 0
high-sensitivity C-reactive protein 391 mg/L | 0
D-dimer >50 000 ng/mL | 0
fibrinogen 439 mg/dL | 0
creatinine kinase myocardial band 31.8 ng/mL | 0
troponin I 0.61 ng/mL | 0
electrocardiogram showed sinus tachycardia | 0
chest X-ray revealed heterogenous consolidation | 0
blood culture | 0
high-flow nasal oxygen therapy | 0
oxygen saturation improved to 92% | 0
respiratory rate improved to 26 breaths per minute | 0
blood pressure improved to 130/80 mmHg | 0
heart rate improved to 120 beats per minute | 0
aspirin therapy | 0
clopidogrel therapy | 0
intravenous unfractionated heparin therapy | 0
activated partial thromboplastin time monitoring | 0
transfer to intensive care unit | 0
meropenem therapy | 0
levofloxacin therapy | 0
dexamethasone therapy | 0
famotidine therapy | 0
vitamin D therapy | 0
ascorbic acid therapy | 0
zinc therapy | 0
atorvastatin therapy | 0
N-acetyl cysteine therapy | 0
nebulized lidocaine therapy | 0
oxygen supplementation down-titrated | 144
simple face mask at 6 liters/minute | 144
blood gas analysis | 144
pH 7.41 | 144
pCO2 37 mmHg | 144
pO2 74 mmHg | 144
HCO3 24 mmol/L | 144
base deficit -1 mmol/L | 144
lactic acid 1.36 mmol/L | 144
procalcitonin decreased to 7.4 ng/mL | 144
high-sensitivity C-reactive protein decreased to 0.13 mg/dL | 144
D-dimer decreased to 5308 ng/mL | 144
fibrinogen increased to 523 mg/dL | 144
alanine aminotransferase decreased to 153 U/L | 144
aspartate aminotransferase decreased to 62 U/L | 144
sudden clinical deterioration | 144
labored breathing | 144
desaturation | 144
hypotension | 144
altered mental status | 144
endotracheal intubation | 144
inotropic and vasopressor agents | 144
computed tomography-pulmonary angiography | 168
thrombosis in bilateral pulmonary arteries | 168
thrombosis in multiple branches of pulmonary veins | 168
brain CT scan | 168
infarct on the cortical-subcortical left parietal lobe | 168
infarct on the pons | 168
infarct on the left part of the cerebellum | 168
rescue thrombolytic therapy with streptokinase | 168
high-sensitivity C-reactive protein increased to 221.1 mg/dL | 336
ferritin >15,000 μg/L | 336
D-dimer decreased to 2597 ng/mL | 336
fibrinogen increased to 634 mg/dL | 336
tocilizumab therapy | 336
death due to multiple end-organ failure | 432