76 years old | 0  
    male | 0  
    hypertension | 0  
    type two diabetes | 0  
    smoking | 0  
    alcoholism | 0  
    fatigue | -720  
    anorexia | -720  
    dyspnea | -720  
    presented to community emergency department | 0  
    temperature 37.8 degrees Celsius | 0  
    heart rate 56 beats per minute | 0  
    blood pressure 132/53 mmHg | 0  
    respiratory rate 40 per minute | 0  
    oxygen saturation 94% on room air | 0  
    bilateral pulmonary crackles | 0  
    white blood cell count 35,000/μL | 0  
    creatinine 1.38 mg/dL | 0  
    troponin-I 0.128 ug/L | 0  
    chest x-ray showed pulmonary edema | 0  
    electrocardiogram showed first degree AV block | 0  
    left bundle branch block | 0  
    no previous for comparison | 0  
    two sets of blood cultures drawn | 0  
    treated with ceftriaxone | 0  
    treated with furosemide | 0  
    supplemental oxygen | 0  
    developed worsening dyspnea | 24  
    third degree heart block | 24  
    transvenous pacing | 24  
    echocardiography demonstrated aortic valve endocarditis | 24  
    transferred to coronary care unit at tertiary care center | 24  
    transesophageal echocardiography confirmed native aortic valve endocarditis | 168  
    vegetation | 168  
    abscess involving non-coronary sinus | 168  
    lateral aspect of the annulus with fistula into left ventricular outflow tract | 168  
    small shunt into the right atrium | 168  
    involvement of mitral-aortic continuity | 168  
    large vegetation extending into left atrium | 168  
    gram negative rods identified in blood cultures | 120  
    MALDI-TOF mass spectrometry identified Capnocytophaga canimorsus | 144  
    sensitive to ceftriaxone | 144  
    sensitive to ampicillin | 144  
    sensitive to ciprofloxacin | 144  
    asked about dog exposure | 144  
    reported repeat severe dog bites over past three months | 144  
    extensive valvular involvement | 0  
    underwent cardiac surgery on post-admission day 10 | 240  
    aortic valve replacement | 240  
    mitral valve repair | 240  
    closure of Sinus of Valsalva aneurysm | 240  
    pathology of aortic valve demonstrated two aortic valve cusps | 240  
    tan-brown confluent vegetations (2.3 cm) | 240  
    cusp perforation (0.8 cm) | 240  
    cusp aneurysm (0.9×0.9×0.8 cm) | 240  
    gram-stain negative | 240  
    bacterial culture of aortic valve negative | 240  
    post-operative blood cultures negative | 240  
    post-operative course uncomplicated | 240  
    discharged on post-admission day twenty | 480  
    planned duration of antimicrobial treatment six weeks | 480  