72 years old | 0
retired mechanic | 0
left shoulder remote rotator cuff injury | 0
adhesive capsulitis | 0
aneurysmal dilation of the ascending aorta | 0
mild aortic insufficiency | 0
crush injury to the left forearm and hand | -96
rib fractures | -96
pneumohemothorax | -96
acute treatment of injuries | -96
transferred to home hospital | -96
admitted to intensive care unit | -96
symptoms of sepsis | -96
left upper extremity infection | -96
preoperative x-ray | -96
plate and screw fixation | -96
significant debris | -96
bone fragments | -96
soft tissue swelling | -96
postoperative day 5 | -48
second surgery | -48
extensive debridement | -48
lavage for deep infection | -48
flexor carpi radialis nonviable | -48
hand intrinsic muscles nonviable | -48
long flexors nonviable | -48
extensors nonviable | -48
wound packed | -48
discussion of limb salvage | -48
transradial amputation discussion | -48
postoperative day 7 | -24
transradial below-elbow amputation | -24
postoperative day 19 | 120
debridement of amputation site | 120
split-thickness skin grafting | 120
discharge home | 120
referral for prosthetic fitting | 120
rehabilitation impaired by PLP | 120
intense sensation of flexion | 120
cramping of digits 1 to 3 | 120
trials of medication | 0
nonpharmacological management | 0
socket modifications | 0
desensitization therapy | 0
compressive stump covers | 0
mirror therapy | 0
discontinuation of prosthesis use | 0
gabapentin titrated to 600 mg three times daily | 0
severe lightheadedness | 0
pregabalin titrated to 150 mg twice daily | 0
tramadol 37.5 mg as needed | 0
hydromorphone 1 mg to 2 mg every 4 h as needed | 0
local xylocaine injections | 0
x-ray of residual limb | 24
heterotopic ossification identified | 24
calcitonin trial | 24
intranasal calcitonin 200 units daily | 24
significant reduction in PLP | 168
discontinued analgesic medication | 168
three-month follow-up | 2160
minimal pain | 2160
no HO progression | 2160
six-month follow-up | 4320
return to prosthesis use | 4320
18-month follow-up | 12960
minimal phantom pain | 12960
continued prosthesis use | 12960
no surgical management | 12960
