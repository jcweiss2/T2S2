55 years old | 0
male | 0
admitted to the hospital | 0
previous history of resection of a right adrenal tumor | -8760
resection of a right adrenal tumor | -8760
post-traumatic hematuria | -8760
mass (diameter 10.6 cm) | -8760
normal blood pressure | -8760
stage II tumor | -8760
follow-up | -8760
annual basis | -8760
computed tomography | -8760
positron emission tomography (PET) | -8760
asymptomatic | -8760
liver enzymes disturbances | -24
abdomen computed tomography | -24
magnetic resonance imaging | -24
large (14.4 × 12.6 cm) intrahepatic mass | -24
no other localization | -24
PET-scan (FDG-18) | -24
metabolically active | -24
liver biopsy | -24
molecular research assay | -24
Tumor Hotspot MASTR Plus | -24
negative | -24
surgical resection of the intrahepatic tumor | 0
pre-anesthetic visit | 0
asymptomatic | 0
normal arterial blood pressure | 0
normal heart rate | 0
no medication | 0
induction of anesthesia | 0
sevoflurane | 0
mobilization of the right liver | 0
severe adhesions | 0
bleeding | 0
hypotensive | 0
blood transfusions | 0
norepinephrine infusion | 0
parenchymal transection | 0
easy | 0
bleeding free | 0
no portal nor hepatic vein was opened | 0
no residual bleeding | 0
cristalloids | 0
colloids | 0
no changes in oxygen saturation | 0
no changes in end-tidal carbon dioxide | 0
no air embolism | 0
intensive care unit (ICU) | 0
norepinephrine infusion rate | 0
arterial blood pressure | 0
fluid replacement therapy | 0
hemoglobin concentration | 0
total plasma protein concentration | 0
refractory vasoplegic shock | 0
transthoracic echocardiography | 0
well preserved left ventricular function | 0
low filling pressures | 0
fluids | 0
vasopressors | 0
methylprednisolone | 0
ventilated | 0
generalized oedema | 24
anuric renal failure | 24
lactic acidosis | 24
four-limb ischemia | 24
rhabdomyolysis | 24
abdominal compartment syndrome (ACS) | 24
bladder pressure | 24
multiple organ dysfunction | 24
second laparotomy | 48
decompression of ACS | 48
no acute liver failure | 48
no intestinal ischemia | 48
blood cultures | 168
Escherichia coli | 168
septic shock | 168
acute respiratory distress syndrome | 168
death | 216
catecholamines | -24
cortisol | -24
synaptophysin + | -24
MART1 + | -24
alpha-inhibin + | -24
CKAE1/AE3 - | -24
chromogranin - | -24
Ki67 index | -24
metastatic adrenocortical carcinoma | -24
postmortem examination | 216
acute tubular necrosis | 216
centrilobular liver necrosis | 216
hemorrhagic necrosis of the spleen | 216
lung congestion | 216
diffuse intra-alveolar hemorrhage | 216
inflammatory cell infiltration | 216
coronary arteries | 216
no signs of inflammatory or ischemic injury | 216
myocardium | 216