28 years old | 0
female | 0
farmer | 0
admitted to the Department of Critical Care Medicine | 0
fever | -168
shortness of breath | -168
spontaneous abortion | -168
IVF-ET treatment | -98
pregnancy established | -98
vaginal bleeding | -9
spontaneous abortion | -7
uterine clearance | -7
feeling cold | -7
chills | -7
cough | -7
dizziness | -7
general fatigue | -7
body temperature 38.7 °C | -7
cefopodoxime proxetil treatment | -7
no improvement | -5
worsening shortness of breath | -2
admitted to local hospital | -1
chest CT scan | -1
scattered ground-glass dense opacities | -1
nodular shadows | -1
referred to emergency department | 0
severe pneumonia diagnosis | 0
anti-infection therapy | 0
oxygen supply | 0
infection-related indices increased | 0
cefoperazone sodium/sulbactam sodium and moxifloxacin treatment | 0
worsening shortness of breath | 0
non-invasive ventilator | 0
dyspnea | 6
irritability | 6
oxygen saturation 44% | 6
arterial blood gas analysis | 6
type I respiratory failure | 6
physical examination | 0
body temperature 36.9 °C | 0
heart rate 123 beats/min | 0
respiratory rate 26 breaths/min | 0
blood pressure 86/54 mmHg | 0
emaciated body | 0
ventilation via ventilator and tracheal tube intubation | 0
rough breathing sound | 0
wet rales | 0
no abnormality in heart and abdominal examination | 0
pitting edema in lower limbs | 0
laboratory test results | 0
imaging results | 0
bedside chest X-ray scan | 0
double-lung pneumonia | 0
fiberoptic bronchoscopy | 0
yellow sputum scabbing | 0
alveolar lavage fluid collection | 0
body temperature 38 °C | 24
noradrenaline treatment | 24
oxygen concentration 80% | 24
sedation and analgesic treatments | 24
PCT increased | 24
CRP level 142.4 mg/L | 24
anti-infection treatment with meropenem and linezolid | 48
improvement in infection indices | 72
PCT 2.24 ng/mL | 72
blood leukocyte count 4.49×10^9/L | 72
neutrophils 82.2% | 72
blood pressure 110/70 mmHg | 72
heart rate 86 bpm | 72
respiration rate 18 breaths/min | 72
SpO2 98% | 72
ventilator use reduced | 72
PEEP 8 cm H2O | 72
FiO2 45% | 72
arterial blood gas analysis | 72
pH 7.438 | 72
PCO2 40.1 mmHg | 72
PO2 118 mmHg | 72
HCO3- 26.8 mmol/L | 72
BE 2.7 mmol/L | 72
lactate 2.0 mmol/L | 72
discharged from ventilator | 72
exercise | 72
fever | 72
CRP 90.5 mg/L | 72
abdominal ultrasonography | 72
pelvic ultrasonography | 72
gynecological ultrasonography | 72
no obvious abnormalities | 72
mNGS test | 72
M. tuberculosis complex group | 72
Xpert results positive | 72
pulmonary TB diagnosis | 72
hematogenous disseminated pulmonary TB | 72
anti-TB therapy | 72
isoniazid | 72
rifampicin | 72
pyrazinamide | 72
ethambutol | 72
chest radiographs | 120
extensive exudation | 120
small nodules | 120
referred to specialized TB hospital | 120
M. tuberculosis culture positive | 120
quadruple anti-TB therapy | 120
ventilator assistance | 120
death | 168
multiple organ failure | 168