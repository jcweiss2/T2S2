38 years old | 0 | 0 
male | 0 | 0 
admitted to the hospital | 0 | 0 
HBV-associated PAN | -156 | 0 
acute abdomen | 0 | 0 
septic shock | 0 | 0 
prednisolone | -4320 | -120 
cyclophosphamide | -4320 | -120 
Tenofovir | -4320 | -168 
chronic renal failure | -156 | 0 
diabetes mellitus Type II | -156 | 0 
free sub diaphragmatic air | 0 | 0 
peritonitis | 0 | 0 
three perforations of the small intestine | 0 | 0 
segmental enterectomy with anastomosis | 0 | 24 
mechanical ventilation | 0 | 72 
circulatory support | 0 | 72 
acute-on-chronic renal failure | 0 | 72 
weaned off the ventilator | 72 | 72 
haemodynamically stable | 72 | 120 
tenofovir orally | 72 | 168 
IV methylprednisolone | 72 | 120 
enteric content from abdominal drain catheter | 168 | 168 
second explorative laparotomy | 168 | 168 
two new perforations | 168 | 168 
multiple areas of patchy necrosis | 168 | 168 
plasma exchanges | 168 | 360 
IV cyclophosphamide | 168 | 168 
IV methylprednisolone | 168 | 192 
IV prednisone | 192 | 360 
third laparotomy | 216 | 216 
three new necrotic lesions | 216 | 216 
necrotic lesion on the left lobe of the liver | 216 | 216 
fourth laparotomy | 264 | 264 
segmental enterectomy with anastomosis | 264 | 264 
cholecystectomy | 264 | 264 
anastomotic leak | 264 | 264 
gangrenous gallbladder | 264 | 264 
septic shock | 360 | 360 
multiple organ failure | 360 | 360 
death | 360 | 360 
weight loss | -8760 | -156 
myalgias | -8760 | -156 
fever | -8760 | -156 
skin erythema | -8760 | -156 
deterioration of renal function | -8760 | -156 
new onset of diabetes mellitus Type II | -8760 | -156 
hypertension | -8760 | -156 
HBsAg | -156 | 0 
HBeAg | -156 | 0 
Anti-HBcAb | -156 | 0 
absence of Anti-HBsAb | -156 | 0 
absence of Anti-HBeAb | -156 | 0