19 years old | 0
female | 0
admitted to the hospital | 0
impaired consciousness | 0
social drinker | -672
frequent diarrhea | -672
abdominal pain | -672
diarrheal symptom worsened | -144
high fever | -72
headache | -72
myalgia | -72
unstable vital signs | 0
blood pressure 70/40 mm Hg | 0
pulse rate 130 beats/min | 0
body temperature 41.0℃ | 0
respiratory rate 35/min | 0
stuporous mental status | 0
diffusely tender and distended abdomen | 0
white blood cell count 21,440/mm3 | 0
neutrophil 92% | 0
hemoglobin 13.4 g/dL | 0
platelet 332,000/µL | 0
urea 10 mg/dL | 0
creatinine 1.1 mg/dL | 0
C-reactive protein 92.9 mg/L | 0
elevated cardiac troponin I | 0
elevated creatine kinase-MB | 0
negative human immunodeficiency virus antibody | 0
negative hepatitis B surface antigen | 0
negative hepatitis C virus antibody | 0
negative anti-nuclear antibody | 0
normal blood and urine cultures | 0
normal stool examinations | 0
sinus tachycardia | 0
interstitial pulmonary edema | 0
dilated ventricles with akinesia | 0
severely impaired systolic function | 0
estimated ejection fraction 38% | 0
fulminant myocarditis with acute LV failure | 0
active inflammatory wall thickening in the distal ileum | 0
associated mesenteric hyperemia | 0
intervening normal segments of the ileum | 0
intubation | 0
ventilator care | 0
intravenous hydration | 0
inotropic support with dopamine | 0
inotropic support with noradrenaline | 0
inotropic support with dobutamine | 0
clinical condition improved | 24
intubation tube removed | 24
decreased cardiac troponin I | 24
viral antibody titers checked | 24
low positive coxsackie virus A4 antibody titer | 24
low positive coxsackie virus A16 antibody titer | 24
low positive coxsackie virus B1 antibody titer | 24
low positive coxsackie virus B3 antibody titer | 24
high positive coxsackie virus B4 antibody titer | 24
low positive adenovirus antibody titer | 24
improved LV systolic function | 168
estimated ejection fraction 62% | 168
discharged | 240
angiotensin-converting enzyme inhibitors | 240
colonoscopy | 672
ulceration with stenosis in the terminal ileum | 672
multiple aphthous ulcers in the rectum | 672
non-caseating granulomatous inflammation | 672
Crohn's disease diagnosis | 672
oral steroids | 672
mesalazine | 672
improved symptoms | 672
maintenance therapy with mesalazine | 672
maintenance therapy with azathioprine | 672
unchanged coxsackie virus B4 antibody titer | 864