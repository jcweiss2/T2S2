70 years old | 0
male | 0
persistent cough | -2160
never smoked | 0
taking statin | -87600
taking anti-hypertensive drugs | -87600
vital signs stable | 0
physical examination no significant findings | 0
chest CT scan | 0
PET scan | 0
malignant lung mass 4.8 cm x 4.3 cm in left lower lobe | 0
multiple mediastinal lymph nodes | 0
bone metastases | 0
stage IV cancer | 0
bronchoscopy irregular mucosal changes | 0
protruding mass at LLL orifice | 0
invasive mucinous lung adenocarcinoma | 0
TTF-1 positive | 0
no EGFR mutations | 0
no ALK fusions | 0
no ROS1 fusions | 0
PD-L1 TPS 100% | 0
first-line pembrolizumab monotherapy initiated | 0
slight increase in primary tumor mass | 264
slight increase in mediastinal lymph nodes | 264
two additional cycles of pembrolizumab | 264
cough difficult to control | 264
antitussives use | 264
inhaled bronchodilators use | 264
systemic corticosteroids use | 264
marked enlargement of primary lung tumor | 528
marked enlargement of mediastinal lymph nodes | 528
newly developed bone metastases | 528
carcinoembryonic antigen elevated to 57.2 ng/mL | 528
frontline treatment discontinued | 528
switched to pemetrexed and carboplatin | 528
NGS performed | 528
KRAS p.G12V mutation | 528
TP53 p.E286K mutation | 528
STK11 p.Y36fs* mutation | 528
pneumonia developed | 528
serum CRP elevated | 528
procalcitonin elevated | 528
bronchial obstruction at LLL | 528
no ground-glass opacities | 528
no airspace consolidations in right lung | 528
intensive care with antibiotics | 528
mechanical ventilation | 528
sepsis | 528
patient succumbed | 528
