58 years old | 0
female | 0
diabetic | 0
admitted to intensive care unit | 0
emergency coronary angiogram | -48
normal coronaries | -48
urinary tract infection | -48
diabetic ketoacidosis | -48
treated for urinary tract infection and diabetic ketoacidosis | -48
pulseless ventricular tachycardia | -48
advanced cardiac life support protocol | -48
transferred for coronary angiogram | -48
troponin levels raised | 0
2D echocardiography showing left ventricular hypokinesia | 0
mechanically ventilated | 0
vasopressors | 0
norepinephrine | 0
easily arousable to call | 0
no neurological deficit | 0
episodes of ill-sustained ventricular tachycardia | 0
arterial blood gas | 0
optimal oxygenation | 0
high anion gap acidosis | 0
neutrophilic leukocytosis | 0
intravenous amiodarone infusion | 0
correction of electrolyte disturbances | 0
hypokalemia | 0
hypomagnesemia | 0
intravenous meropenem | 0
human insulin infusion | 0
controlling blood sugar levels | 0
general condition improved | 12
resolution of shock | 12
correction of acidosis | 12
restoration of normal sinus rhythm | 12
extubated | 12
computed tomography urography | 12
pyelonephritis | 12
bedside 2D echocardiography | 12
Takotsubo cardiomyopathy | 12
apical ballooning of the left ventricle | 12
speckle tracking on echocardiography | 12
apical hypokinesia | 12
electrophysiologist opinion | 12
oral bisoprolol | 12
oral amiodarone | 12
shifted to step-down unit | 24
cardiac magnetic resonance imaging | 24
Takotsubo cardiomyopathy appearance | 24
mid and apical cavity | 24
shifted back to intensive care unit | 36
episodes of ill-sustained ventricular tachycardia | 36
synchronized cardioversion | 36
intravenous antiarrhythmic bolus doses | 36
amiodarone | 36
lignocaine | 36
thoracic epidural catheter | 36
sympathetic blockade | 36
ropivacaine | 36
hypokalemia | 36
no further episodes of ventricular tachycardia | 84
Holter monitoring | 84
epidural catheter removed | 108
discharged from hospital | 216
oral propefenone | 216
amiodarone | 216
bisoprolol | 216
two dimensional echocardiography | 216
mild apical and distal interventricular septal hypokinesia | 216
ejection fraction 45% | 216