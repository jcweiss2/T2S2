67 years old | 0
male | 0
hypertension | -672
degenerative joint disease | -672
bilateral knee replacement | -672
substance abuse | -672
trauma to his face and chest wall | -24
lightheadedness | 0
fatigue | 0
leukocytosis | 0
hemoglobin of 10.2 g | 0
venous lactic acid of 2.4 mol/l | 0
intramuscular and subpectoral hematoma | 0
extrapleural extension into the chest | 0
acute right second through fifth anterior rib fractures | 0
bilateral lower lobe bronchopneumonia | 0
blood cultures | 0
intravenous piperacillin–tazobactam | 0
afebrile | 0
hypotensive | 0
admitted to the intensive care unit | 0
suspected septic shock | 0
initiation of vasopressors | 0
intravenous vancomycin | 48
cefepime | 48
metronidazole | 48
repeat blood cultures | 48
repeat urine cultures | 48
repeat sputum cultures | 48
methicillin-resistant Staphylococcus aureus | 48
intravenous vancomycin | 96
left knee pain | 120
notable swelling on physical exam | 120
sterile left knee aspiration | 120
synovial fluid cloudy | 120
amber colored | 120
white blood cells of 9.28 × 103/mcL | 120
6.0 × 103/mcL | 120
calcium pyrophosphate crystals | 120
complete washout and debridement of the joint | 144
retention of the prosthesis | 144
infected knee | 144
purulence | 144
intravenous cefazolin | 168
C. bifermentans | 240
intravenous ampicillin–sulbactam | 240
oral suppression with amoxicillin–clavulanic acid | 240
contrast computerized tomography scan of the abdomen | 240
human immunodeficiency virus screening | 240
discharged to a rehabilitation facility | 384
full range of motion of his left knee | 1056
no signs of lingering joint or systemic infection | 1056
taking Augmentin | 1056
medication adherence | 1056