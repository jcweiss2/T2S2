40 years old | 0
female | 0
admitted to the hospital | 0
DLBCL | -720
R-CHOP treatment | -720
fever | -4320
high fever | -4320
shortness of breath | 0
moist rales | 0
body temperature 37.8 ℃ | 0
blood pressure 162/104 mmHg | 0
pulse 147 bpm | 0
respiratory rate 28 breaths/min | 0
white blood cell count 7.17 × 10^9/L | 0
red blood cell count 2.86 × 10^12/L | 0
haemoglobin level 95 g/L | 0
platelet count 403 × 10^9/L | 0
C-reactive protein level 277.6 mg/L | 0
bone marrow cytology | 0
lymphoid malignant tumour cells 22.5% | 0
CD20 (+) | 0
TDT (-) | 0
anti-infective treatment | 0
imipenem 1 g q6h+ | 0
tigecycline 100 mg q12h+ | 0
carprofen 5 mg qd | 0
body temperature 36.5 °C | 24
oxygen saturation 91.3% | 24
white blood cell count 12.32 × 10^9/L | 24
lymphocyte classification 1.0% | 24
monocyte classification 1.0% | 24
neutrophil classification 97.0% | 24
CRP level 79.0 mg/L | 24
Pneumocystis jirovecii | 0
Legionella pneumophila | 0
coinfection | 0
septic shock | 168
drug-induced pancreatitis | 168
enlarged pancreas | 168
echo changes | 168
endotracheal intubation ventilator | 24
discharged | -720
death | 720
Pneumocystis pneumonia | 0
Legionella infection | 0
next-generation sequencing | 0
metagenomic next-generation sequencing | 0
Illumina NextSeq 550 | 0
SE75 sequencing strategy | 0
pathogenic microorganism database | 0
informed consent | -720
Research Ethics Committee | -720