60 years old | 0
lady | 0
presented to the emergency department | 0
migratory right lower quadrant pain | -24
diarrhea | -24
fevers | -24
rigors | -24
previous diverticulitis | 0
hypertension | 0
shocked | 0
blood pressure of 86/52 | 0
borderline tachycardiac at 95 bpm | 0
tender in the right lower quadrant | 0
guarding | 0
acute kidney injury (AKI) | 0
eGFR of 37 ml/min | 0
white cell count of 32.9 (109/L) | 0
referred to the surgical team | 0
clinical diagnosis of acute appendicitis | 0
Alvarado score of nine | 0
urine microscopy showed >500 leucocytes | 0
non-contrast computer tomography (CT) performed | 0
malrotated right ectopic kidney | 0
perinephric stranding | 0
non-obstructing 6 mm calculus in renal pelvis | 0
treated with ampicillin | 0
reduced dose of gentamicin | 0
persisting shock | 0
admitted to the intensive care unit (ICU) | 0
inotropic support | 0
urine culture grew Escherichia coli | 0
blood culture grew Escherichia coli | 0
repeat CT with contrast performed | 0
persisting high fevers | 0
severe right lower quadrant pain | 0
early renal abscess | 0
ongoing sepsis | 0
absence of urology service | 0
transferred to another hospital | 0
insertion of a ureteric stent | 0
continued to improve post stent insertion | 0
discharged when clinically well | 0
removal of stone | 1008
ureteric stent 6 weeks later | 1008
