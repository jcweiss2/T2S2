43 years old | 0
male | 0
admitted to the hospital | 0
fever | 0
ascites | 0
sickle cell anemia | -9360
splenectomy | -9360
cholecystectomy | -9360
transit ischemic attack | -7920
diagnostic imaging control with CT scan | 0
giant mass in the left upper-abdominal quadrant | 0
CT-angio with i.v. contrast infusion | 0
giant splenic aneurysm | 0
concomitant contrast infusion into the enlarged splenic vein | 0
diagnostic centesis | 0
aspirin treatment | -24
hydroxyurea treatment | -24
tazobactam treatment | -24
omeprazole treatment | -24
spironolactone treatment | -24
rifaximin treatment | -24
saccharomyces boulardii treatment | -24
enoxaparin treatment | -24
surgery | 24
open repair via supra-infraumbilical incision | 24
intraperitoneal access to the aorta | 24
covered rupture | 24
4 liters of ascites and blood in the peritoneal cavity | 24
sac preparation | 24
omentum and aneurysmatic sac removal | 24
cross clamp to the orifice of the splenic artery | 24
vessels ligation | 24
post-operative care in ICU | 48
transfer to General Surgery Department | 72
portal vein thrombosis | 72
antithrombotic treatment modification | 72
transfer to Internal Medicine Department | 240
fever | 312
high levels of laboratory inflammation markers | 312
paralytic ileus | 312
low Hct | 312
diagnostic imaging control with CT and DSA | 312
minor signs of bleeding in the area of the stomach atrium | 312
hemorrhagic pancreatitis | 312
investigative laparotomy | 312
intraperitoneal lavage | 312
VAC of the abdominal cave | 312
transfer to ICU | 312
sepsis treatment | 432
transfer to General Surgery Department | 672
discharge | 720