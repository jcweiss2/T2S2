32 years old | 0
male | 0
Vietnamese | 0
admitted to the hospital | 0
abdominal pain | 0
syncope | 0
hypotension | 0
systolic blood pressure 50+ | 0
smoker | -8760
2-pack year history | -8760
occasional drinker | -8760
technician in a factory | -8760
severely tender and tense abdomen | 0
free fluid | 0
large 8x9cm AAA | 0
CT aortogram | 0
tortuous and aneurysmal dilatation of the abdominal aorta | 0
10.8 × 10.8 cm in axial dimension | 0
24.1 cm in cranio-caudal length | 0
extending into the left common iliac artery | 0
involving the origin of the bilateral renal arteries | 0
large retroperitoneal hematoma | 0
emergency open abdominal aortic aneurysm repair | 0
aortic cross clamp | 0
bifurcated aortic graft | 0
anastomosed proximally | 0
distally to the bilateral common iliac arteries | 0
on table angiogram of the left lower limb | 0
abrupt cut-off at the level of the left popliteal artery | 0
transverse arteriotomy | 0
Fogarty balloon catheter | 0
multiple thrombi | 0
final angiogram | 0
in-line flow to the foot via the anterior tibial artery | 0
foot pulses were palpable and strong | 0
transferred to the intensive care unit | 0
extubated on post-operative day 1 | 24
intensive chest physiotherapy | 24
incentive spirometry | 24
nasogastric feeding on POD2 | 48
oral diet by POD 6 | 144
fever | 96
piperacillin-tazobactam | 96
negative septic work up | 120
down-trending inflammatory markers | 120
pro-calcitonin level within normal limits | 120
surgical sites were healing well | 120
no hematoma or signs of infection | 120
acute kidney injury | 0
managed with proper hydration | 0
normalising of his renal function | 0
transient liver enzyme rise | 0
resolved gradually | 0
coagulation profile was preserved | 0
clinically stable | 288
independently mobile | 288
fit for discharge from hospital | 288
discharged | 288
histopathological examination | 288
degenerative changes of the aortic wall | 288
consistent with aortic rupture | 288
no granulomas | 288
no giant cells | 288
no obliterative phlebitis | 288
no storiform fibrosis | 288
no malignancy | 288
no evidence of any infective process | 288
multiple investigations | 0
lost to follow up | 288
genetic testing | 288
pectus excavatum | 0
arachnodactyly | 0
pes planus | 0
keloid at the midline laparotomy wound | 288
elevated C-reactive protein | 0
elevated erythrocyte sedimentation rate | 0
normal serum cholesterol | 0
normal homocysteine level | 0
no evidence of atheroma | 0
no tell-tale clinical features of rheumatological disorders | 0
no vasculitis | 0
no dry eyes | 0
no xerostomia | 0
no abnormal hair loss | 0
no rashes | 0