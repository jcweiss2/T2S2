52 years old | 0
male | 0
admitted to the hospital | 0
watery diarrhea | -96
chills | -96
fever | -96
eating slices of raw fish | -96
drinking soju | -6720
cefotaxime | -48
fever persisted | -48
blisters | -48
referred to the hospital | -24
admitted to the ICU | 0
body temperature of 38°C | 0
blood pressure of 73/40 mmHg | 0
pulse rate of 100 beats per minute | 0
respiratory rate of 40 breaths /min | 0
mild pallor | 0
icteric sclera | 0
blisters with ecchymosis | 0
hematocrit level of 26.6% | 0
white blood cell count of 3,230 cells/mm3 | 0
platelet count of 41,000 cells/mm3 | 0
pH of 7.306 | 0
carbon dioxide tension of 25.7 mmHg | 0
partial pressure of oxygen of 29.7 mmHg | 0
bicarbonate level of 13.0 mmol/L | 0
base excess of 11.4 mmol/L | 0
oxygen saturation level of 49.7% | 0
lactic acid level of 15.8 mmol/L | 0
C-reactive protein concentration of 6.52 mg/dL | 0
procalcitonin concentration of 57.030 ng/mL | 0
total bilirubin of 2.85 mg/dL | 0
direct bilirubin of 2.3 mg/dL | 0
alkaline phosphatase of 65 U/dL | 0
aspartate transaminase of 181 U/dL | 0
alanine transaminase of 35 U/dL | 0
albumin of 2.5 g/dL | 0
total protein of 5.6 g/dL | 0
prothrombin time of 25.1 s | 0
partial thromboplastin time of 85.5 s | 0
international normalize ratio of 2.32 | 0
urea nitrogen of 34.4 mg/dL | 0
creatinine of 3.66 mg/dL | 0
hemoglobin A1c of 5.2% | 0
newly formed pulmonary shadows | 6
intravenous corticosteroid therapy | 0
inotropic agents | 0
empirical intravenous antibiotic therapy | 0
cefepime | 0
doxycycline | 0
metabolic acidosis | 12
arterial blood gas analysis | 12
pH of 7.388 | 12
carbon dioxide tension of 23.5 mmHg | 12
bicarbonate level of 14.3 mmol/L | 12
oxygen saturation level of 83.8% | 12
ventilator therapy | 12
tracheal intubation | 12
blood pressure restored | 24
hemorrhagic blisters | 24
continuous renal replacement therapy | 24
metabolic acidosis worsened | 48
multiple organ failure | 48
arterial blood gas analysis | 48
pH of 7.100 | 48
carbon dioxide tension of 40.9 mmHg | 48
partial pressure of oxygen of 71.6 mmHg | 48
bicarbonate level of 12.4 mmol/L | 48
base excess of 17.2 mmol/L | 48
oxygen saturation level of 88.1% | 48
lactic acid level of 19.5 mmol/L | 48
aspartate aminotransferase of 5,852 U/dL | 48
alanine aminotransferase of 455 U/dL | 48
total bilirubin of 7.22 mg/dL | 48
direct bilirubin of 5.65 mg/dL | 48
creatine phosphokinase of 75,885 U/L | 48
lactate dehydrogenase of 8,433 U/L | 48
died of septic shock | 72
V. cholerae non-O1/O139 infection | 0
Gram-negative rods | 0
VITEK II Compact | 0
serological tests | 0
polymerase chain reaction test | 0
cholera toxin gene | 0
V. cholerae O139 O antigen-specific gene | 0
V. cholerae O1 O antigen-specific gene | 0
Daegu Public Health and Environment Research Institute | 0