74 years old | 0  
    woman | 0  
    admitted to the Intensive Care Unit | 0  
    severe respiratory dysfunction | 0  
    diffuse alveolar infiltrates | 0  
    dyspnea on exertion | -1464  
    dry cough | -48  
    chest pain | -48  
    myalgias | -8760  
    malaise | -8760  
    anorexia | -8760  
    polymyalgia rheumatica | -8760  
    prednisolone | -8760  
    tachypneic | 0  
    central cyanosis | 0  
    use of inspiratory accessory muscles | 0  
    bilateral inspiratory crackles | 0  
    severe hypoxemia | 0  
    pH 7.48 | 0  
    partial pressure of oxygen 49 mmHg | 0  
    partial pressure of carbon dioxide 31 mmHg | 0  
    oxygen saturation 83% | 0  
    anemia | 0  
    hemoglobin level 10.9 g/dL | 0  
    leukocytosis | 0  
    white blood cell count 11.5x10^9/L | 0  
    normal platelet count 213x10^9/L | 0  
    elevated erythrocyte sedimentation rate 80 mm/h | 0  
    elevated C-reactive protein 3710 mg/dL | 0  
    impaired kidney function | 0  
    serum creatinine 1.73 mg/dL | 0  
    diffuse bilateral patchy opacities | 0  
    normal sinus radiographs | 0  
    admitted to Pulmonary Department | 0  
    severe lower respiratory tract infection | 0  
    intravenous ceftriaxone | 0  
    intravenous azithromycin | 0  
    worsening respiratory insufficiency | 0  
    noninvasive ventilation | 0  
    high-resolution computed tomography | 0  
    ground-glass opacities | 0  
    consolidation in right upper lobe | 0  
    subpleural sparing | 0  
    normal abdomen computed tomography | 0  
    clinical condition deteriorated | 96  
    transferred to ICU | 96  
    worsening respiratory distress | 96  
    commencing circulatory failure | 96  
    APACHE II score 24 | 0  
    intubated | 96  
    mechanical ventilation | 96  
    pressure control ventilation 22 cm H2O | 96  
    positive end-expiratory pressure 8 | 96  
    PaO2/FiO2 125 | 96  
    ARDS | 96  
    cardiovascular support | 96  
    fluids | 96  
    vasopressors | 96  
    significant decline of hemoglobin 7.9 g/dL | 96  
    marked leukocytosis | 96  
    white blood cell count 18.5x10^9/L | 96  
    worsening renal function | 96  
    creatinine 2.06 mg/dL | 96  
    active urine sediment | 96  
    dysmorphic red blood cells | 96  
    red blood casts | 96  
    negative transthoracic echocardiogram | 96  
    normal left ventricular systolic function | 96  
    clinical stabilization | 96  
    fiberoptic bronchoscopy | 96  
    no endobronchial lesions | 96  
    hemorrhagic bronchoalveolar lavage fluid | 96  
    negative bacterial cultures | 96  
    negative mycobacterial cultures | 96  
    no cytological evidence of malignancy | 96  
    blood in stool | 96  
    colonoscopy | 96  
    gut biopsy | 96  
    mild edema | 96  
    histopathologic changes of chronic colitis | 96  
    ANCA positive PR3-cANCA | 96  
    titer 1/80 | 96  
    negative antiglomerular basement membrane | 96  
    negative antinuclear antibodies | 96  
    negative extractable nuclear antigens | 96  
    negative hepatitis B serology | 96  
    negative hepatitis C serology | 96  
    rheumatoid factor 10 IU/mL | 96  
    normal complement levels | 96  
    diagnosed with ANCA-associated vasculitis | 96  
    pulmonary-renal syndrome | 96  
    high-dose steroids | 96  
    intravenous methylprednisolone | 96  
    prednisone | 96  
    cyclophosphamide | 96  
    plasmapheresis | 96  
    clinical stabilization | 240  
    improvement of arterial blood gases | 240  
    resolution of ARDS | 240  
    weaned from mechanical ventilation | 240  
    referred to rehabilitation unit | 960  
    died of sepsis | 960  
    nosocomial pneumonia | 960  
    no hospital discharge | 960  
    