47 years old | 0
female | 0
admitted to the hospital | 0
weakness | -7
numbness of the limbs | -7
nausea | -7
fatigue | -7
dyspnea | -7
fever | -7
cough | -7
diagnosed with acute upper respiratory infection | -7
influenza virus A | -7
history of GBS | -2520
GBS caused by influenza virus A | -2520
clear consciousness | 0
blood pressure 84/58 mmHg | 0
heart rate 115 beats/minute | 0
peripheral oxygen saturation 99% | 0
respiratory rate 22 breaths/minute | 0
body temperature 35.7°C | 0
manual muscle testing revealed strength of 3/5 in both lower extremities | 0
manual muscle testing revealed strength of 4/5 in both upper extremities | 0
electrocardiogram revealed sinus tachycardia | 0
elevated ST segment in lead V2-6 | 0
cardiothoracic ratio 53% | 0
pulmonary congestion | 0
high levels of troponin I | 0
high levels of brain natriuretic peptides | 0
elevated creatine kinase | 0
elevated creatine kinase-myocardial band | 0
positive influenza virus A | 0
fulminant myocarditis | 0
venoarterial extracorporeal membrane oxygenation | 0
intra-aortic balloon pumping | 0
sedation | 0
norepinephrine | 0
severely reduced LV function | 6
ejection fraction of 4% | 6
liver enzyme level increased | 72
bilirubin increased | 72
aspartate aminotransferase increased | 72
alanine aminotransferase increased | 72
improved | 120
left ventricular ejection fraction of 67% | 120
weaned from VA-ECMO | 168
weaned from IABP | 168
weaned from ventilator | 264
motor and sensory disorders in her limbs remained | 192
manual muscle testing revealed further reduced muscle strength | 192
absent deep tendon reflexes | 192
sensory disturbance was glove-and-stocking type | 192
nerve conduction study revealed decreased amplitude | 192
axonal GBS | 192
immunoadsorption for GBS | 216
motor and sensory disorders gradually improved | 216
discharged | 648