papillary thyroid carcinoma | -9840 | -9840 | Factual
resection | -9840 | -9840 | Factual
radiotherapy | -9840 | -9840 | Factual
stenosis of the esophagus | -6720 | 0 | Factual
repeated aspiration | -6720 | 0 | Factual
respiratory insufficiency | -6720 | 0 | Factual
pneumonia | -6720 | 0 | Factual
purulent pleurisy | -6720 | 0 | Factual
pleurectomy | -6720 | 0 | Factual
restrictive ventilation pattern | -6720 | 0 | Factual
recurrent nerve palsy | -6720 | 0 | Factual
percutaneous endoscopic gastrostomy | -6720 | -6720 | Factual
tracheostoma | -6720 | -6720 | Factual
home ventilation | -6720 | 0 | Factual
decreased mobility | -4380 | 0 | Factual
secondary depression | -4380 | 0 | Factual
stented left axis vertebralis | -2190 | -2190 | Factual
stenosis of the internal axis carotis | -2190 | 0 | Factual
arterial hypertension | -2190 | 0 | Factual
secondary lactase deficiency | -2190 | 0 | Factual
esophageal stenosis dilation | -168 | -168 | Factual
decreasing general condition | 0 | 0 | Factual
fistula between the esophagus and tracheal membrane | 0 | 0 | Factual
pneumonia by 4-multiresistente gramnegative Pseudomonas aeruginosa | 0 | 0 | Factual
veno-venous extracorporeal membrane oxygenation | 0 | 720 | Factual
ventilation through a tracheostoma | 0 | 720 | Factual
thoracic computed tomography | 24 | 24 | Factual
big fistula of the tracheal membrane | 24 | 24 | Factual
endobronchial stenting | 48 | 48 | Factual
retrograde stenting | 48 | 48 | Factual
Freitag stent placement | 48 | 48 | Factual
regular tracheal cannula introduction | 72 | 72 | Factual
spontaneous breathing work increase | 120 | 600 | Factual
vv-ECMO support reduction | 120 | 600 | Factual
lungs re-aerated | 120 | 600 | Factual
patient woke up | 120 | 600 | Factual
communication with family | 120 | 600 | Factual
infections continued | 120 | 720 | Factual
spontaneous work of breathing never exceeded 170 mL per breath | 120 | 720 | Factual
reduction of intravenous saline injection | 600 | 720 | Factual
vv-ECMO support reduction | 600 | 720 | Factual
patient died | 720 | 720 | Factual
pulmonary infection | 720 | 720 | Factual