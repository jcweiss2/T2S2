62 years old | 0
female | 0
Ph + ALL | -2160
bone marrow biopsy | -2160
flow cytometry | -2160
induction chemotherapy | -2160
hyper-CVAD | -2160
vincristine | -2160
doxorubicin | -2160
dexamethasone | -2160
intrathecal methotrexate | -2160
nonoliguric acute kidney injury | -672
discontinued hyper-CVAD | -672
oral dasatinib | -672
continued intrathecal methotrexate | -672
headaches | -48
neck pain | -48
back pain | -48
low-grade fever | -48
worsening generalized weakness | -48
increased difficulty with ambulation | -48
confusion | -48
last dose of intrathecal methotrexate | -96
febrile | 0
tachycardic | 0
normotensive | 0
diaphoretic | 0
lethargic | 0
neck stiffness | 0
hemoglobin 6.9 g/dL | 0
transfused with one unit of packed red blood cells | 0
white blood cell count 6.8 K/uL | 0
computed tomography imaging | 0
no acute process | 0
contraindication of having an implanted spinal stimulator | 0
started on cefepime | 0
started on vancomycin | 0
started on ampicillin | 0
prophylactic fluconazole | 0
prophylactic acyclovir | 0
attempted lumbar puncture | 24
confused | 24
unable to cooperate with the procedure | 24
transferred to ICU | 24
agitated | 24
required rapid sequence intubation | 24
mechanical ventilation | 24
lumbar puncture | 48
cerebrospinal fluid cultures showed no growth | 48
negative PCR for herpes simplex virus | 48
negative PCR for varicella-zoster virus | 48
negative PCR for Lyme disease | 48
negative PCR for West Nile virus | 48
negative upper respiratory panel | 48
negative influenza testing | 48
negative SARS-CoV-2 PCR | 48
gradually improved | 120
remained hemodynamically stable | 120
discontinued antimicrobial therapy | 120
extubation | 120
transitioned from ICU to general ward | 216
encephalopathic | 216
mentation rapidly improved | 216
profoundly physically weak | 216
nasogastric tube removed | 240
began to tolerate an oral diet | 240
physical and occupational therapy | 240
able to stand up with assistance | 264
no confusion or agitation | 288
back to baseline mentation | 288
fever resolved | 288
leukocytosis resolved | 288
recommended for rehabilitation therapy | 288
declined rehabilitation therapy | 288
provided with home health care | 288
no further episodes of encephalopathy | 720
ceased intrathecal methotrexate | 720
maintained on dasatinib | 720
started on blinatumomab | 720