47 years old | 0
female | 0
multiparous | 0
menorrhagia | -672
adenomyosis | -672
total laparoscopic hysterectomy | -672
bilateral salphingoopherectomy | -672
watery leakage per vaginally | -48
cystoscopy | -48
trigonal vesicovaginal fistula | -48
patulous right ureteric orifice | -48
transvaginal VVF repair | -48
Martius flap interposition | -48
discharged | -336
catheter | -336
static cystogram | 0
right loin pain | 336
fever | 336
chills | 336
urosepsis | 336
readmitted | 336
resuscitated | 336
blood culture | 336
urine culture | 336
Escherichia Coli | 336
retrospective inspection | 336
plain X-ray | 336
Foley's catheter | 336
dilated right ureter | 336
contrast extravasation | 336
subcapsular region | 336
right kidney | 336
deflated | 336
repositioned | 336
fluoroscopic guidance | 336
plain computed tomography | 336
CT KUB | 336
curvilinear right subcapsular collection | 336
perinephric stranding | 336
absence of periureteric extravasation | 336
intravenous antibiotics | 336
intensive care unit | 336
recovered | 720
discharged | 720
voiding well | 720
no leakage of urine | 720