63 years old | 0
male | 0
admitted to the hospital | 0
hypertension | -6720
chronic back pain | -6720
spinal stenosis | -6720
lower extremity edema | -6720
oxycodone | -6720
losartan | -6720
furosemide | -840
fever | -336
diffuse maculopapular rash | -168
cough | -168
profuse watery diarrhea | -336
hematochezia | -336
abdominal pain | -336
dry nonproductive cough | -168
fevers up to 38.6°C | -168
stopped taking furosemide | -168
temperature of 38.6°C | 0
blood pressure 126/59 mm Hg | 0
heart rate 103 beats per minute | 0
respiratory rate 22 breaths per minute | 0
oxygen saturation was 95% | 0
diffuse erythematous maculopapular rash | 0
tachycardia | 0
leukocytosis of 11.8×10^9/L | 0
elevated eosinophil count of 1.29×10^9/L | 0
hemoglobin and platelets were normal | 0
creatinine, electrolyte, and liver enzymes tests were all normal | 0
inflammatory markers were elevated | 0
C-reactive protein (CRP) of 229 | 0
erythrocyte sedimentation rate (ESR) of 31 | 0
blood gas showed hypoxemia | 0
partial oxygen was 66 mm Hg | 0
computed tomography (CT) scan of the chest showed significant hilar lymphadenopathy | 0
interstitial changes consistent with pneumonitis | 0
levofloxacin | 0
intravenous (IV) fluids | 0
doxycycline | 24
skin biopsy | 24
thrombocytopenia | 24
atrial fibrillation with rapid ventricular response | 48
re-exposure to furosemide | 48
worsening rash | 60
worsening hypoxia | 60
increased fever | 60
increased eosinophil count | 60
increased creatinine | 60
acute kidney injury | 60
DRESS syndrome secondary to furosemide | 120
oral prednisone 1 mg/kg daily | 120
discharged | 360
atovaquone | 360
spironolactone | 360
improved symptomatically | 1008
laboratory testing normalized | 1008
fatigue | 1008
mild shortness of breath | 1008
insomnia from steroids | 1008