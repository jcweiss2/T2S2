67 years old | 0
    man | 0
    admitted to the hospital | 0
    mucosal resection for early gastric cancer | -10080
    partial resection for left lung cancer | -10080
    collected knee-high wild grass from a riverbed for 10 days | -672
    systemic pain | -504
    fatigue | -504
    fever | -336
    chills | -336
    watery diarrhea | -336
    loss of appetite | -336
    mildly disturbed consciousness | -336
    visited the department of internal medicine | -168
    decreased white blood cells (WBC) | 0
    platelet counts | 0
    elevated hepatic enzyme levels | 0
    hepatic dysfunction | 0
    hospitalized | 0
    height of 169.0 cm | 0
    body weight of 52.3 kg | 0
    Glasgow Coma Scale of 14: E3, V5, M6 | 0
    blood pressure of 130/79 mmHg | 0
    heart rate (HR) of 96/min | 0
    regular pulse | 0
    respiratory rate (RR) of 20/min | 0
    O2 saturation (SPO2) of 94% in room air | 0
    temperature of 38.9°C | 0
    no remarkable head-and-neck abnormalities | 0
    no chest abnormalities | 0
    crusted skin lesions on the medial surface of the left thigh | 0
    freely movable adenopathy of approximately 2 cm in size without tenderness | 0
    aggregated papules in the right inguinal region | 0
    no remarkable neurological abnormalities | 0
    blood count: 1,300 /μL WBC | 0
    platelets: 30,000 /μL | 0
    neutrophil count: 899 /μL | 0
    lymphocyte count: 342 /μL | 0
    activated partial thromboplastin time (APTT) of 48.2 seconds | 0
    mild increase in C-reactive protein (CRP) levels at 1.3 mg/dL | 0
    elevated aspartate aminotransferase (AST) at 230 U/L | 0
    elevated lactate dehydrogenase (LDH) at 760 U/L | 0
    elevated creatine kinase (CK) at 746 U/L | 0
    chest radiography normal | 0
    electrocardiography normal | 0
    simple head-and-neck computed tomography (CT) scan normal | 0
    suspected sepsis | 24
    suspected febrile neutropenia (FN) | 24
    associated with hemophagocytosis | 24
    administered antibiotics | 24
    elevated ferritin levels of 15,165 ng/mL | 48
    screened for antibodies specific for cytomegalovirus | 48
    screened for antibodies specific for Epstein-Barr virus (EBV) | 48
    blood culture negative | 48
    bone marrow biopsy performed | 48
    hemophagocytosis | 48
    fewer mature myeloid series cells | 48
    more monocytoid cells | 48
    more lymphoid cells | 48
    immunohistological examination revealed CD3- and CD4-positive T cells | 48
    MUM-1-positive lymphoid cells | 48
    CD68-positive histiomonocytes | 48
    CD163-positive histiomonocytes | 48
    no EBV-encoded small RNAs (EBERs)-positive cells detected | 48
    diagnosed with HLH | 48
    administered prednisolone (PSL) at 60 mg/day | 48
    gradually tapered PSL | 72
    stopped PSL on day 12 of administration | 288
    developed chest pain | 72
    shivering | 72
    fever of 39.2°C | 72
    blood pressure at 88/52 mmHg | 72
    HR at 89/min | 72
    RR at 24/min | 72
    SPO2 at 94% (6-L mask for oxygen administration) | 72
    elevated CK levels at 953 U/L | 72
    elevated LDH at 1,405 U/L | 72
    high-sensitivity troponin I (TnI) at 271 pg/mL | 72
    transthoracic echocardiography showed severe left ventricular dysfunction (LVEF of 15%) | 72
    electrocardiogram (ECG) showed slight ST elevation in V1-2 leads | 72
    contrast-enhanced CT of chest and abdomen normal | 72
    fulfilled diagnostic criteria of clinically suspected myocarditis | 72
    acute myocarditis suspected | 72
    did not perform coronary angiography (CAG) | 72
    did not perform EMB | 72
    continued respiratory and circulatory management | 72
    continued infection control in ICU | 72
    TnI peaked at 82.6 pg/mL | 72
    suspected SFTS | 72
    submitted serum, urine samples, and throat swabs to public health center | 72
    moved to negative-pressure room | 72
    RT-PCR detected 1.77×106 SFTSV RNA copies/mL | 72
    submitted bone marrow sections to National Institute of Infectious Disease | 72
    infected cells stained positively by anti-SFTSV-nucleoprotein (N) antibody | 72
    considered steroid pulse therapy for HLH with SFTS | 72
    did not proceed with steroid pulse therapy | 72
    withdrew from circulatory agonist | 336
    withdrew from ventilator management | 336
    ECG improvement of ST elevation in V1-2 leads | 336
    submitted serum confirmed negativity for viremia | 408
    released from quarantine | 408
    performed CAG | 576
    performed EMB | 576
    no coronary artery stenosis observed | 576
    myocardium mildly hypertrophic | 576
    mild myofibrillar loss | 576
    mild myofibrillar disarrangement | 576
    no active mononuclear cell infiltration adjacent to damaged myocardium | 576
    immunohistochemistry revealed increases in CD3-positive T cells (10/mm2) | 576
    increases in CD68-positive macrophages (18/mm2) | 576
    tenascin-C expression in stroma | 576
    myocardial tissues immunostaining negative for anti-SFTSV antibody | 576
    discharged | 696
    follow-up transthoracic echocardiography showed EF of 52.5% | 1176
    no heart failure thereafter | 1176
    <|eot_id|>
    