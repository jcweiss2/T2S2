22 years old | 0
female | 0
Malay ethnicity | 0
admitted to the haematology department | 0
fever | -168
left axillary swelling | -168
no past medical history | 0
no family history | 0
non-smoker | 0
does not consume alcohol | 0
works as a bank clerk | 0
pale | 0
left axillary swelling of 5 x 5 cm | 0
firm | 0
non-tender | 0
no discharge | 0
no palpable lymph nodes | 0
no organomegaly | 0
normochromic normocytic anaemia | 0
leucocytosis | 0
thrombocytopenia | 0
no coagulopathy | 0
blasts in peripheral blood smear | 0
abnormal promyelocytes in peripheral blood smear | 0
faggot cells in peripheral blood smear | 0
blasts in bone marrow aspirate | 0
abnormal promyelocytes in bone marrow aspirate | 0
faggot cells in bone marrow aspirate | 0
hypercellular marrow | 0
blast population expressing myeloperoxidase | 0
lacking CD34 | 0
lacking CD3 | 0
cluster of aberrant myeloid cells expressing CD117 | 0
cluster of aberrant myeloid cells expressing cMPO | 0
cluster of aberrant myeloid cells expressing CD13 | 0
cluster of aberrant myeloid cells expressing CD33 | 0
cluster of aberrant myeloid cells expressing CD38 | 0
lacking CD34 | 0
lacking HL-DR | 0
PML-RAR-alpha fusion gene | 0
t(15;17) (q22; q12) | 0
diffuse monomorphic infiltrates | 0
neoplastic cells exhibiting fine nuclear chromatin | 0
moderate rim of basophilic cytoplasm | 0
positive for MPO | 0
positive for CD13 | 0
positive for CD33 | 0
positive for CD68 | 0
positive for CD117 | 0
negative for CD34 | 0
negative for HLA-DR | 0
granulocytic sarcoma | 0
high-risk APML | 0
diagnosed with high-risk APML | 0
treated with dexamethasone | 0
treated with all-trans-retinoic-acid | 0
treated with arsenic trioxide | 0
treated with idarubicin | 0
developed culture-negative neutropenic sepsis | 336
Type 1 respiratory failure | 336
intubated | 336
nursed at the intensive care unit | 336
no evidence of alveolar haemorrhage | 336
diffuse nodular pulmonary infiltrations | 336
no features of pulmonary embolism | 336
serum galactomannan not detected | 336
treated with antimicrobials | 336
responded completely to antimicrobials | 336
completed induction therapy | 720
completed consolidation therapy | 1000
completed maintenance therapy | 2000
in complete molecular remission | 2000
in complete molecular remission for 2 years | 2000