61 years old | 0
    male | 0
    bipolar disorder | -43800
    lithium carbonate medication (600 mg/day) | -43800
    Emergency Unit admission | 0
    progressively decreased consciousness level | -120
    lithium overdose | 0
    sleepiness | -48
    prostration | -48
    mental confusion | -48
    rigidity of the lower extremities | -48
    insulin therapy | -43800
    metformin 850 mg 3xday | -43800
    thyroxine (T4) 50 mcg/day | -43800
    enalapril 40 mg/day | -43800
    atenolol 100 mg/day | -43800
    non-pale | 0
    anicteric | 0
    acyanotic | 0
    rales in pulmonary base | 0
    respiratory rate 29 bpm | 0
    irregular cardiac rhythm | 0
    heart rate 130 bpm | 0
    blood pressure 80/40 mmHg | 0
    hemoglobin 12.5 g/dL | 0
    hematocrit 36% | 0
    WBC 9500/mm³ | 0
    neutrophils 82% | 0
    lymphocytes 18% | 0
    platelets 207,000/mm³ | 0
    negative blood cultures | 0
    normal chest X-radiography | 0
    lithium poisoning | 0
    hemodialysis | 24
    lithium serum level 2.9 mmol/L | 24
    creatinine 2.3 mg/dL | 24
    urea 114 mg/dL | 24
    potassium 3.1 mEq/L | 24
    sodium 145 mEq/L | 24
    mechanical ventilation | 24
    dopamine administration | 24
    hypotension | 24
    bradycardia | 24
    normal brain tomography | 24
    metabolic encephalopathy | 24
    echocardiogram showing dilated left atrium and left ventricular hypertrophy | 24
    normal left ventricular systolic function | 24
    CKMB 132 U/L | 24
    cardiac troponin I 20.92 μg/L | 24
    cardiac catheterization | 24
    normal coronary circulation | 24
    ECG atrial fibrillation | 0
    ST segment elevation 1 mm diffusely | 0
    T-wave inversion | 0
    left ventricular overload | 0
    atrial fibrillation with low-ventricular response | 24
    bradycardia 45 bpm | 24
    tachycardia 174 bpm | 24
    electrical cardioversion | 24
    ventricular tachycardia | 72
    bradyarrhythmia | 72
    temporary pacemaker implantation | 72
    pacemaker turned off | 96
    serum lithium levels 0.6 mmol/L | 96
    sinus rhythm | 96
    absence of arrhythmias | 96
    tracheostomy | 96
    hemorrhagic complications | 120
    cardiorespiratory arrest | 120
    pulseless electrical activity | 120
    unsuccessful resuscitation | 120
    death | 120

<|eot_id|>