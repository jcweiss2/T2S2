62 years old | 0
female | 0
ulcerative colitis | 0
5E-ASA | 0
acute severe flare of UC | -672
infliximab | -672
CT findings | -672
positive serology for pANCA | 0
positive serology for ANA | 0
breast carcinoma | 0
family history of UC | 0
fever | 0
cough | 0
vomiting | 0
diarrhea | 0
generalized weakness | 0
confusion | 0
lethargy | 0
low GCS score (12/15) | 0
acutely altered mental status | 0
mild neck stiffness | 0
baseline bloods | 0
chest X-ray | 0
septic screen | 0
blood cultures | 0
urine cultures | 0
elevated CRP (94 mg/dL) | 0
stable hemoglobin (12.8 g/dL) | 0
COVID-19 not detected | 0
lower respiratory tract infection | 0
intravenous piperacillin/tazobactam | 0
fluids | 0
new-onset confusion | 0
persistent hypotension | 0
admitted to ICU | 0
blood cultures positive for L. monocytogenes | 0
brain CT | 0
no acute intracranial pathology | 0
lumbar puncture | 0
cloudy cerebrospinal fluid | 0
elevated WBC count (1,600/mm3) | 0
CSF glucose (1.8 mmol/L) | 0
CSF protein (1.75 g/L) | 0
bacterial meningitis | 0
L. monocytogenes DNA detected | 0
flare of colitis | 720
Mayo 3 endoscopic appearance | 720
L. monocytogenes sepsis | 0
meningeal involvement | 0
infliximab held | 0
intravenous amoxicillin | 0
discontinued infliximab | 0
recovered from meningitis | 0
vedolizumab commenced | 720
discussion of colectomy | 720
acute flare of severe UC | 1440
Mayo 3 on endoscopy | 1440
subtotal colectomy | 1440
unremarkable post-surgical course | 1440
