71 years old | 0 | 0 
female | 0 | 0 
admitted to the hospital | 0 | 0 
unconscious state | 0 | 0 
history of hypertension | 0 | 0 
history of ischaemic heart disease | 0 | 0 
history of peripheral vascular disease | 0 | 0 
stroke | 0 | 0 
head computed tomographic scan | 0 | 0 
condition deteriorated | 48 | 48 
inotropic support | 48 | 48 
septic shock | 48 | 48 
elevated levels of inflammatory markers | 48 | 48 
erythrocyte sedimentation rate | 48 | 48 
C-reactive protein | 48 | 48 
blood culture | 48 | 48 
yeast in blood culture | 48 | 48 
caspofungin | 48 | 72 
died | 72 | 72 
Lodderomyces elongisporus | 48 | 72 
identification by VITEK 2 yeast identification system | 48 | 72 
identification by CHROMagar Candida | 72 | 72 
identification by acetate ascospore agar | 72 | 72 
identification by PCR sequencing of ITS region of rDNA | 72 | 72 
antifungal susceptibility | 72 | 72 
amphotericin B | 72 | 72 
fluconazole | 72 | 72 
voriconazole | 72 | 72 
posaconazole | 72 | 72 
itraconazole | 72 | 72 
flucytosine | 72 | 72 
caspofungin | 72 | 72 
micafungin | 72 | 72 
hospitalization for lower limb ischaemia | -336 | -336 
discharge from hospital | -168 | -168 
history of heart disease | 0 | 0 
history of stroke | 0 | 0 
no antibiotics | 0 | 72 
no central lines | 0 | 72 
fungaemia | 48 | 72 
inoculation of yeast from skin | -72 | 48 
translocation from gastrointestinal tract | -72 | 48 
endocarditis | 0 | 0 
global prevalence | 0 | 0 
isolation from patients in distant geographic regions | 0 | 0 
turquoise blue colonies on CHROMagar Candida | 72 | 72 
ellipsoidal to elongate ascospores on acetate ascospore agar | 72 | 72 
Candida parapsilosis complex | 0 | 0 
reduced susceptibility to echinocandins | 0 | 0 
in vitro MIC values | 72 | 72 
antifungal therapy | 48 | 72 
outcome | 72 | 72 
mortality rates | 72 | 72 
diagnostic challenges | 0 | 0 
therapeutic challenges | 0 | 0 
delay in accurate identification | 0 | 0 
lack of experience in management | 0 | 0 
prophylactic use of antifungal agents | 0 | 0 
therapeutic use of antifungal agents | 48 | 72 
selection pressure | 0 | 0 
increased colonization | 0 | 0 
invasive infection | 48 | 72 
rare yeast infections | 0 | 0 
higher mortality rates | 72 | 72 
technical support | 0 | 0 
Mycology Reference laboratory | 0 | 0 
S. Varghese | 0 | 0 
S. Vayalil | 0 | 0 
O. Al-Musallam | 0 | 0