65 years old | 0
male | 0
hypertension | 0
COPD | 0
Parkinson's disease | 0
irregular treatment | 0
follow-up | 0
respiratory distress | -168
productive cough | -168
hypercapnic respiratory failure | 0
altered sensorium | 0
leukocytosis | 0
intubated | 0
invasive mechanical ventilation | 0
ventilator-associated pneumonia | 216
Acinetobacter baumanii | 216
cefoperazone/sulbactam | 216
colistin | 216
fall in procalcitonin levels | 216
spontaneous breath trial (SBT) failed | 216
worsening respiratory acidosis | 216
desaturation | 216
hypotension | 216
hypovolemic hypotension | 216
polyuria | 216
hypokalemia | 216
hyponatremia | 216
hypocalcemia | 216
hypomagnesaemia | 216
high fractional excretion of sodium (FeNa) | 216
transtubular potassium gradient (TTKG) | 216
excess renal loss of electrolytes | 216
parenteral correction of electrolytes | 216
recurrence | 216
stopping colistin | 216
parameters started to reverse | 240
extubated | 240
grade III bed sores | 240
infected | 240
Klebsiella spp. | 240
sepsis | 648
rising procalcitonin levels | 648
restarted on colistin | 648
electrolyte abnormalities | 648
polyuria | 648
hypovolemic hypotension | 648
supraventricular tachycardia (SVT) | 648
low level of serum magnesium | 648
magnesium replacement | 648
no recurrence | 648
course of 10 day colistin | 648
repeated electrolyte corrections | 648
volume replacements | 648
discharged | 1008
resolution of abnormalities | 1008