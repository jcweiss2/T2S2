abruptio placenta | -168
emergency cesarean delivery | -168
birth | 0
Apgar 4 | 0
Apgar 8 | 5
respiratory distress | 0
CPAP | 0
respiratory distress syndrome | 0
ground-glass opacity | 0
minor respiratory acidosis | 0
surfactant | 0
bowel movement | 12
trophic feeding | 72
abdominal distension | 144
tachycardia | 144
tachypnea | 144
thrombocytopenia | 144
neutropenia | 144
C-reactive protein 70 mg/L | 144
meropenem | 144
vancomycin | 144
antibiotics discontinued | 216
feeding restarted | 216
high-flow oxygen | 336
unexplained apnea | 504
unexplained apnea | 672
septic examination negative | 504
septic examination negative | 672
brain MRI normal | 504
nasogastric tube | 504
conjugated hyperbilirubinemia | 504
neonatal cholestasis workup | 504
hepatitis and total parenteral nutrition suspected | 504
genetic studies | 504
X-ray of spine normal | 504
echocardiogram normal | 504
eye test normal | 504
skull X-ray craniosynostosis | 504
hepatosplenomegaly not seen | 504
biliary atresia not seen | 504
albumin level decline | 504
bilirubin rise | 504
AST rise | 504
ALT rise | 504
albumin infusions | 504
ursodeoxycholic acid | 504
infectious etiology investigation | 504
TSH normal | 504
T3 normal | 504
T4 normal | 504
cortisol normal | 504
metabolic disorders negative | 504
galactosemia negative | 504
tyrosinemia type 1 negative | 504
whole-exome sequencing | 1008
severe cyanosis | 1176
apnea | 1176
bradycardia | 1176
cardio-respiratory resuscitation | 1176
intubation | 1176
mechanical breathing | 1176
epinephrine | 1176
septic shock | 1176
multiorgan failure | 1176
disseminated intravascular coagulation | 1176
acute renal damage | 1176
capillary leak syndrome | 1176
death | 2400
whole-exome sequencing results | 2407
NOTCH2 gene mutation | 2407
heterozygous variant c.1076c>T | 2407
Ser359Phe | 2407
chr1: 120512166 | 2407
ALGS2 diagnosis | 2407