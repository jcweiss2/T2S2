12 years old | 0
neutered female | 0
American cocker spaniel | 0
presented for evaluation | 0
dyspnea | -48
anorexia | -48
gallbladder mucocele | -192
pancreatitis | -192
extrahepatic bile duct obstruction | -192
gallbladder mucocele surgically removed | -168
discharged | -96
lethargic | 0
tachypnea | 0
respiratory distress | 0
heart rate 128 bpm | 0
heart murmur not auscultated | 0
SpO2 not measurable | 0
systolic blood pressure 162 mmHg | 0
diastolic blood pressure 69 mmHg | 0
leukocytosis 38.3 × 103/µl | 0
thrombocytopenia 103 × 103/µl | 0
serum biochemical profile within normal range | 0
prothrombin time 8.0 sec | 0
activated partial thromboplastin time 21.1 sec | 0
fibrinogen 344 mg/dl | 0
thoracic radiographs revealed cardiac enlargement | 0
enlargement of main pulmonary artery | 0
interstitial and alveolar lung patterns | 0
transthoracic echocardiography performed | 0
severe RV dilation | 0
right atrial dilation | 0
main pulmonary artery dilation | 0
RV to left ventricular end-diastolic basal diameter ratio 1.17 | 0
myocardial hypokinesis of RV free wall | 0
interventricular septal flattening | 0
paradoxical septal motion | 0
mild tricuspid regurgitation | 0
TR velocity 4.6 m/sec | 0
RA pressure estimated 10 mmHg | 0
systolic PA pressure estimated 93.4 mmHg | 0
PA acceleration time 35 msec | 0
PA ejection time 204 msec | 0
acceleration time/ejection time ratio 0.17 | 0
mitral regurgitation not identified | 0
transmitral flow pattern impaired relaxation | 0
RV function indices impaired | 0
RV-SD increased | 0
CT angiography performed | 0
filling defect in left and right main PA | 0
filling defect in brachiocephalic veins | 0
atelectasis in middle lobe | 0
ground-grass opacity in lung lobes | 0
diagnosed as acute PTE | 0
severe pulmonary hypertension | 0
treated in intensive care unit | 0
oxygen therapy initiated | 0
low molecular heparin administered | 0
cefazolin administered | 0
aspirin administered | 0
clopidogrel administered | 0
respiratory status improved | 216
good clinical condition on day 9 | 216
breathing normally in room air | 216
echocardiographic variables improved | 216
reduction in right heart size | 216
improvement in interventricular septal flattening | 216
TR velocity decreased to 2.9 m/sec | 216
hypokinesis of RV free wall improved | 216
RV dyssynchrony improved | 216
CT angiography on day 9 | 216
filling defects unchanged | 216
lung field abnormalities resolved | 216
discharged on day 10 | 240
plasma D-dimer elevated 7.19 µg/ml | 0
fibrin degradation product elevated 24.0 µg/ml | 0
acute PTE after surgery and prolonged cage rest | 0
