4 years old | 0
    intact male | 0
    Golden retriever | 0
    weight 32 kg | 0
    admitted to a local animal hospital | 0
    abdominal distention | -168
    melena | -168
    lethargy | -168
    anorexia | -168
    raised indoors | -168
    no toxicant exposure | -168
    azotemia | -168
    hypoalbuminemia | -168
    administration of 6% hydroxyethyl starch 130/0.4 solution | -168
    increased creatinine level | -168
    proteinuria | -168
    azotemia persisted | -168
    proteinuria persisted | -168
    referred to Veterinary Medical Teaching Hospital | 336
    severe azotemia | 336
    ascites | 336
    gastrointestinal bleeding | 336
    normothermic (38.0°C) | 336
    normal heart rate (120 bpm) | 336
    normal respiratory rate (30/min) | 336
    hypertensive (175 mmHg) | 336
    ecchymosis | 336
    distended abdomen | 336
    microcytic non-regenerative anemia | 336
    neutrophilia | 336
    thrombocytopenia | 336
    hypoalbuminemia | 336
    hypoproteinemia | 336
    hyperbilirubinemia | 336
    increased alkaline phosphatase | 336
    increased gamma glutamyl transferase | 336
    increased fasting bile acid | 336
    mild increased activated partial thromboplastin | 336
    deteriorated azotemia | 336
    hyperphosphatemia | 336
    metabolic acidosis | 336
    hyponatremia | 336
    hyperkalemia | 336
    hypocalcemia | 336
    hyposthenuria | 336
    proteinuria | 336
    anuria | 336
    increased renal cortex echogenicity | 336
    liver assessment disturbance due to ascites | 336
    ascites removal | 336
    transudate ascites | 336
    chronic liver failure suspected | 336
    decreased functional liver enzymes | 336
    coagulopathy | 336
    globulin within reference interval | 336
    cholesterol within reference interval | 336
    no marked proteinuria on day 2 | 336
    acute anuric renal failure | 336
    decreased liver function | 336
    euthanized | 336
    necropsy performed | 336
    multifocal hepatic nodules | 336
    petechial-to-ecchymotic hemorrhages in heart | 336
    gastrointestinal bleeding | 336
    renal cortex degeneration | 336
    hepatic fibrosis | 336
    hepatic calcium deposits | 336
    renal tubular necrosis | 336
    glomerular injury | 336
    albumin transudation | 336
    osmotic nephrosis lesions | 336
    acute kidney injury confirmed | 336
    liver cirrhosis confirmed | 336
    platelet dysfunction suspected | 336
    HES-induced AKI | 336
    HES administration controversy in veterinary medicine | 336
    no adverse effects evidence in animals | 336
    lower adverse outcome prevalence in animals | 336
    higher serum amylase activity in dogs | 336
    shorter hospital duration in animals | 336
    hypotheses of HES-induced AKI mechanisms | 336
    osmotic nephrosis hypothesis | 336
    reversible osmotic nephrosis lesions | 336
    pathological evidence of HES-induced injury | 336
    platelet dysfunction causes uncertain | 336
    liver cirrhosis influence on AKI | 336
    warning against synthetic colloids in animals with decreased kidney function | 336
    need for HES adverse effects studies in veterinary medicine | 336
    multicentre studies recommended | 336

    <|eot_id|>
    