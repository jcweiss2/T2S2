64 years old | 0
male | 0
admitted to the hospital | 0
cough | -72
chest X-ray findings with right pleural effusion and a right hilar mass | -72
facial edema | -72
SVC syndrome | -72
transbronchial biopsy | -72
diagnosis of SCLC | -72
right hilar, mediastinal, right supraclavicular, aortic, and superior mediastinal lymph node metastasis | -72
pleural effusion | -72
no brain metastases | -72
no abnormal findings in the abdomen | -72
extensive SCLC | -72
carboplatin | 0
etoposide | 0
right pneumothorax | 96
chest tube drainage | 96
fever | 144
right thoracic empyema | 144
ampicillin/sulbactam | 144
febrile neutropenia | 192
meropenem | 192
filgrastim | 192
pleural effusion culture showed a meropenem-sensitive peptostreptococcus infection | 192
diarrhea | 456
fecal culture | 456
Clostridium difficile toxin | 456
CD antigen | 456
bloody stools | 576
abdominal pain | 576
abdominal CT | 576
intestinal retention | 576
intussusception in the ileocecal region | 576
abscess in the left hepatic lobe | 576
emergency surgery | 600
extensive necrosis of the colon | 600
extensive colectomy | 600
colostomy | 600
septic shock | 600
intensive care management | 600
piperacillin/tazobactam | 600
vancomycin | 600
micafungin | 600
portal vein thrombosis | 672
anticoagulation therapy | 672
Entamoeba histolytica trophozoites | 672
severe inflammatory cell infiltration | 672
abscess formation | 672
bleeding | 672
fibrin | 672
loss of continuity of the intestinal wall | 672
no history of amoebiasis | 0
no sexual intercourse with homosexuals, commercial sex workers, or an unspecified number of people | 0
traveled to the Philippines seven years before the onset of symptoms | -5040
traveled to the West Coast of the United States, Hawaii, and Shanghai 10 years previous | -8760
metronidazole | 792
improved general condition | 1008
liver abscess | 1008
percutaneous catheter drainage | 1008
bacterial culture of the right pleural effusion | 1176
chest tube removal | 1176
paromomycin | 1032
anti-cystic therapy | 1032
lower gastrointestinal endoscopy | 1464
mild white mucus | 1464
residual redness | 1464
carcasses of amoebic trophozoites | 1464
improved general condition | 1464
liver abscess shrank | 1464
palliative radiotherapy | 1404
SVC syndrome exacerbated | 1404
second cycle of chemotherapy | 2016
carboplatin | 2016
etoposide | 2016
partial response | 2016
no recurrence of amoebic dysentery | 2016