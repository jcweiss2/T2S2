63 years old | 0
male | 0
admitted to the hospital | 0
abrupt onset of fever | -24
progressive mental obtundation | -24
Glasgow Coma Scale score 4 | 0
right-sided otitis media | 0
purulent discharge | 0
temperature 36.8° C | 0
pulse 124 | 0
respiration 20 | 0
blood pressure 137/79 mmHg | 0
mild divergent strabismus | 0
eye deviation to the left | 0
deep tendon reflexes symmetric and enhanced | 0
Babinski's sign negative | 0
leukocyte count 18.5 × 10^9/L | 0
neutrophils 91% | 0
monocytes 7% | 0
lymphocytes 3% | 0
red blood cell count 4.7 × 10^12/L | 0
hemoglobin 143 g/L | 0
platelets 172 × 10^9/L | 0
erythrocyte sedimentation rate 80 per h | 0
C-reactive protein 75.5 mg/L | 0
fibrinogen 4.13 g/L | 0
prothrombin time normal | 0
partial-thromboplastin time normal | 0
serum lactate 6.0 mmol/L | 0
magnesium 0.5 mmol/L | 0
phosphorus 0.43 mmol/L | 0
total bilirubin normal | 0
aminotransferases normal | 0
lactate dehydrogenase normal | 0
glucose normal | 0
alkaline phosphatase normal | 0
serum protein electrophoresis normal | 0
blood sodium 134 mmol/L | 0
potassium 3.0 mmol/L | 0
chloride 97 mmol/L | 0
urea nitrogen 5.0 mmol/L | 0
creatinine 88 μmol/L | 0
CSF white cells 200,000 per cubic millimeter | 0
CSF polymorphonuclear cells 95% | 0
CSF glucose 0.0 mmol/L | 0
CSF total protein 12.1 g/L | 0
CSF lactate 15.9 mmol/L | 0
intravenous ceftriaxone 4 g per day | 0
intravenous dexamethasone 48 mg/day | 0
penicillin-resistant Streptococcus pneumoniae cultured from CSF | 0
ceftriaxone-sensitive Streptococcus pneumoniae cultured from CSF | 0
native brain CT scan normal | 0
contrast-enhanced brain CT scan normal | 0
transcranial Doppler ultrasonography | 0
absent diastolic blood flow velocities in both MCA | 0
systolic BFV 25 cm/s left MCA | 0
systolic BFV 23 cm/s right MCA | 0
pulsatility index 4.3 left MCA | 0
pulsatility index 3.4 right MCA | 0
