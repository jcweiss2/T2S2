73 years old | 0  
    male | 0  
    presented to a community hospital | 0  
    jaundice | 0  
    mass in the pancreas | 0  
    obstruction of the common bile duct | 0  
    obstruction of the pancreatic duct | 0  
    no signs of metastases | 0  
    endoprosthesis placed endoscopically in the bile duct | 0  
    brush cytology obtained | 0  
    adenocarcinoma | 0  
    developed severe progressive muscle weakness of his legs | 168  
    developed severe progressive muscle weakness of his arms | 168  
    no pain | 168  
    no loss of sensation | 168  
    no skin abnormalities | 168  
    confined to a wheelchair | 168  
    not able to stand | 168  
    not able to walk | 168  
    diabetes mellitus type 2 | -  
    spontaneous subdural hematoma | -  
    surgically drained subdural hematoma | -  
    family history of breast carcinoma | -  
    family history of colon carcinoma | -  
    creatinine kinase level of 12,570 U/l | 0  
    aspartate aminotransferase 594 U/l | 0  
    alanine aminotransferase 523 U/l | 0  
    lactate dehydrogenase 648 U/l | 0  
    C-reactive protein 11 mg/l | 0  
    magnetic resonance imaging showed diffuse edema in upper muscles | 0  
    magnetic resonance imaging showed diffuse edema in lower leg muscles | 0  
    muscle biopsy revealed numerous necrotic fibers infiltrated by macrophages | 0  
    muscle biopsy revealed few lymphocytes | 0  
    regenerating fibers | 0  
    membrane attack complex positive fibers | 0  
    MHV-I positive non-necrotic muscle fiber | 0  
    skin histology revealed no abnormalities | 0  
    excluded dermatomyositis | 0  
    diagnosis of NAM | 0  
    cooccurrence of NAM with cholangiocarcinoma | 0  
    high-dose dexamethasone therapy started | 0  
    prednisone 20 mg per day | 0  
    intravenous immunoglobulin 2 g/kg | 0  
    laparoscopic pancreatoduodenectomy performed | 0  
    R0 resected pT3N0M0 distal cholangiocarcinoma | 0  
    no adjuvant chemotherapy | 0  
    discharged to a rehabilitation center | 240  
    pancreatic fistula | 240  
    percutaneous drain placed | 240  
    drain removed | 672  
    muscular strength slowly increased postoperatively | 672  
    able to walk a few steps | 672  
    pneumonia | 1008  
    treated with antibiotics | 1008  
    confined to a wheelchair again | 1008  
    admitted to intensive care unit | 1344  
    pneumosepsis | 1344  
    enteral tube feeding | 1344  
    no signs of recovery | 1344  
    discontinued all medical treatment | 1344  
    death | 2880  