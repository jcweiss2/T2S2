38 years old | 0
    male | 0
    obese | 0
    BMI 35.93 kg/m2 | 0
    no known medical or surgical history | 0
    presented to hospital | 0
    fever | -48
    dry cough | -48
    shortness of breath | -48
    positive COVID-19 PCR test | 0
    not received immunization against COVID-19 | 0
    vitally stable on examination | 0
    normal chest examination | 0
    normal cardiovascular examination | 0
    no abdominal tenderness | 0
    chest X-ray | 0
    pneumonic consolidation left lower lobe | 0
    respiratory distress | 96
    tachycardia 100 beats per minute | 96
    tachypnea 36 breaths per minute | 96
    hypotension 90/54 mm Hg | 96
    hypoxia 82% oxygen saturation | 96
    bilateral crepitations | 96
    soft lax abdomen | 96
    repeat chest X-ray | 96
    bilateral patchy infiltrates | 96
    severe COVID-19 pneumonia | 96
    worsening clinically | 96
    worsening radiologically | 96
    started enoxaparin 80 mg subcutaneously twice daily | 96
    severe persistent abdominal pain | 120
    abdominal pain not relieved by analgesia | 120
    abdominal pain not relieved by proton pump inhibitors | 120
    diaphoresis | 120
    vomiting | 120
    vitally stable | 120
    GCS 15/15 | 120
    lax abdomen | 120
    mild epigastric tenderness | 120
    D-dimer 12.91 μg/mL | 120
    persistent pain | 120
    urgent abdominal CT-angiogram | 120
    hypodense filling defect superior mesenteric artery | 120
    hypodense filling defect superior mesenteric vein | 120
    arterial thrombosis | 120
    venous thrombosis | 120
    ischemic changes small bowel loops | 120
    exploratory laparotomy | 120
    ischemic nonviable bowel from duodenojejunal flexure to mid transverse colon | 120
    resected ischemic bowel | 120
    transferred to surgical ICU | 120
    postoperative sepsis | 144
    postoperative multiorgan failure | 144
    pulseless ventricular tachycardia | 144
    resuscitation per ACLS | 144
    no return of spontaneous circulation | 144
    patient passed away | 216
    <|eot_id|>
    