33 years old | 0
female | 0
nausea | -24
vomiting | -24
abdominal pain | -24
discharged | -36
hospitalized | -36
recurrent pericarditis | -36
colchicine | -36
febrile | 0
hypotensive | 0
leukocytosis | 0
elevated serum lactate | 0
acute kidney injury | 0
acute transaminitis | 0
severe coagulopathy | 0
normal serum troponin | 0
negative toxicology screen | 0
normal sinus rhythm | 0
normal biventricular function | 0
sepsis suspected | 0
fluid resuscitated | 0
broad-spectrum antibiotics | 0
vasopressor therapy | 0
multisystem organ failure | 24
intubated | 24
paralyzed | 24
intravascular volume repletion | 24
intravenous vasopressors | 24
stress-dose steroids | 24
high-dose vitamin B12 | 24
Swan-Ganz catheter | 24
distributive shock | 24
cardiogenic shock | 48
high filling pressures | 48
low CO | 48
high systemic vascular resistance | 48
elevated troponin | 48
severe biventricular failure | 48
intravenous milrinone | 48
CRRT | 48
PRBC transfusion | 72
improved CO | 96
decreased troponin | 96
improved multisystem organ failure | 96
neutropenic | 120
recovered LVEF | 144
weaned from vasopressors | 312
taken off CRRT | 312
extubated | 312
hair loss | 576
admitted to taking colchicine | 576
elevated serum colchicine | 30
elevated whole blood colchicine | 14
hypertension | 0
pulmonary emboli | 0
polysubstance abuse | 0
recovered | 720