30 years old | 0
female | 0
pregnant | 0
admitted to the Department of Obstetrics and Pregnancy Pathology | 0
nausea | -72
vomiting | -72
abdominal pain | 0
abdominal distension | 0
moderate tenderness | 0
empirical antibiotic therapy with intravenous ceftriaxone | 0
limited ultrasound | 0
full fetal anatomy assessment | 0
dilated loops of the colon and sigmoid colon | 24
fluid-gas levels | 24
tarry stools | 24
gastroscopy | 24
septic shock | 24
antimicrobial and antifungal treatment | 24
surgical consultation | 24
transferred to the general surgery clinic | 24
surgical treatment | 48
midline laparotomy | 48
moderate amount of serous fluid | 48
dilated large intestine | 48
ruptures of the serosal membrane | 48
appendectomy | 48
cecostomy | 48
safety drains | 48
intraoperatively diagnosed with acute intestinal pseudo-obstruction | 48
respiratory insufficiency | 48
transferred to the Intensive Care Unit | 48
intubated and mechanically ventilated | 48
sedation | 48
enteral and parenteral nutrition | 48
antibiotic therapy | 48
improvement in general condition | 72
transferred to the Department of Surgery | 72
transferred to the obstetrics ward of a lower-level referral hospital | 168
delivered a healthy baby | 1344
procedure to restore the continuity of the gastrointestinal tract | 504
released adhesions | 504
discharged | 504
epilepsy | -8760
mild intellectual disability | -8760
hypothyroidism | -8760
surgical treatment for achalasia of the cardia | -720
Heller cardiomyotomy | -720
Dor fundoplication | -720
long-term pharmacological treatment for epilepsy | -8760
valproic acid | -8760
oxcarbazepine | -8760
thyroid hormone supplementation | -8760