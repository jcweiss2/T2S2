71 years old | 0
male | 0
admitted to the hospital | 0
mild abdominal pain | -72
nausea | -72
profuse diarrhea | -72
abdominal pain worsened | -24
diarrhea worsened | -24
unresponsive | -24
hypotensive | 0
tachycardic | 0
severe pain in lower abdomen | 0
tenderness | 0
no fever | 0
no masses | 0
no lymph nodes | 0
metabolic acidosis | 0
serum lactate level over 6 mmol/L | 0
intravenous fluid reanimation | 0
abdominal computed tomography (CT) | 0
bowel dilated | 0
no free liquid | 0
no air | 0
no masses | 0
abdominal pain worsened | 0
abdominal distention worsened | 0
surgical consultation | 0
surgery | 0
intestinal ischemia | 0
laparotomy | 0
small bowel purplish color | 0
small bowel edematous | 0
no perforation | 0
no necrosis | 0
mesentery engorged | 0
ecchymosis | 0
bowel peristalsis | 0
reanimation maneuvers | 0
second-look surgical laparotomy | 0
Bogota bag | 0
low-molecular-weight heparin | 0
transferred to intensive care unit | 0
angio-3D reconstruction | 0
vascular malformation of superior mesenteric artery | 0
celiacomesenteric trunk | 0
no thrombus | 0
no embolus | 0
second laparotomy | 24
bowel loops better condition | 24
bowel regained normal color | 24
bowel regained mobility | 24
ventilator-associated pneumonia | 24
sepsis | 24
refractory shock | 24
organ failure | 24
death | 24