37 years old | 0
female | 0
posterior occipital lesion | -6720
low-grade glioma with pilocytic features | -6720
occipital craniotomy | 0
supratentorial approach | 0
debulking of the tumor | 0
ASA II | 0
physical exam unremarkable | 0
no allergies | 0
left parietal craniotomy | -8760
partial excision of the tumor | -8760
chemotherapy | -8760
radiotherapy | -8760
increase in intracranial pressure | -4080
external ventricular drainage device insertion | -4080
general anesthesia | -4080
no complications | -4080
recurrence of the brain tumor | -240
right occipital craniotomy | -240
sitting position | -240
general anesthesia | -240
no postoperative complications | -240
blurred vision | -120
metastatic sub-thalamic brain tumor | -120
navigation-assisted tumor debulking | 0
occipital craniotomy | 0
sitting position | 0
minimal head flexion | 0
throat pack insertion | 0
invasive monitoring | 0
left radial arterial line | 0
right subclavian central line | 0
propofol | 0
fentanyl | 0
cisatracurium | 0
cuffed ETT | 0
mechanical ventilator | 0
isoflurane | 0
cisatracurium | 0
remifentanil infusion | 0
Ringer lactate | 0
packed red blood cells | 0
stable vital signs | 0
systolic blood pressure | 0
PaCO2 | 0
oxygen saturation | 0
residual muscle paralysis reversed | 0
neostigmine | 0
atropine | 0
throat pack removed | 0
spontaneous breathing | 0
extubation | 0
bedside neurological exam | 0
left-sided weakness | 0
neurosurgery team informed | 0
repositioning of the patient | 0
relieving mechanical pressure | 0
ischemia reperfusion injury | 0
severe upper airway edema | 0
macroglossia | 0
tongue size increase | 0
O2 saturation decrease | 0
manual mask ventilation | 0
foreign body suspected | 0
oropharynx checked | 0
enlarged tongue | 0
edematous soft palate | 0
epiglottis and vocal cords not visible | 0
intubation difficult | 0
mask ventilation harder | 0
inspiratory stridor | 0
O2 saturation drop | 0
help called | 0
urgent tracheostomy | 0
tracheostomy done | 0
transferred to ICU | 24
mechanical ventilation | 24
sedation | 24
propofol | 24
remifentanil | 24
antibiotics | 24
cefuroxime | 24
vancomycin | 24
levofloxacin | 24
dexamethasone | 24
antihistamine | 24
enteral feeding | 24
nasogastric tube | 24
chest physiotherapy | 24
swollen tongue and neck | 48
mouth gag applied | 48
MRA ordered | 48
MRA not done | 48
increase in WBC count | 120
septic work-up | 120
gram negative bacilli | 120
tongue size increase again | 216
ulcerations on the surface | 216
sepsis | 384
multi-organ failure | 384
asystole | 384
death declared | 384