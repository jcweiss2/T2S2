68 years old | 0
female | 0
admitted to the hospital | 0
AML | -672
bone marrow biopsy | -672
white blood cell count 175,000 | -672
peripheral blasts 27% | -672
normal karyotype | -672
positive for DNMT3, NPM1, PTPN11, and two TET2 pathogenic mutations | -672
induction chemotherapy | -672
decitabine | -672
venetoclax | -672
nonsustained ventricular tachycardia | -672
rapid atrial fibrillation | -672
bacterial pneumonia | -672
maculopapular rash | -24
leukemia cutis | -24
monocytic blasts 44% | -24
nonproductive cough | -24
rhinorrhea | -24
sore throat | -24
afebrile | -24
respiratory viral polymerase chain reaction (PCR) panel positive for SARS-CoV-2 | -24
COVID-19 | -24
mRNA-1273 vaccine | -280
admitted to the medicine service | -24
management of COVID-19 | -24
computed tomography of the chest | -24
no definitive findings of pneumonia | -24
remdesivir | -24
transferred to the malignant hematology service | -17
7+3 reinduction chemotherapy | 0
cytarabine | 0
idarubicin | 0
prophylactic intrathecal cytarabine | 28
retested for COVID-19 | 3
sotrovimab | 3
persistent SARS-CoV-2 positivity | 3
chest pain | 7
computed tomography of the chest | 7
pericarditis | 7
colchicine | 7
blood cell counts reached nadir | 9
absolute neutrophil count (ANC) 0 | 9
neutropenic fever | 20
infectious workup | 20
empiric cefepime | 20
antimicrobial prophylaxis | 20
valacyclovir | 20
isavuconazole | 20
levofloxacin | 20
counts started recovering | 25
ANC 170 | 25
infectious control monitored COVID-19 threshold (CT) count | 25
discharged | 36
COVID-19 PCR retested | 36
recovery bone marrow biopsy | 36
morphologic complete remission | 36
persistent mutations involving DNMT3 and TET2 | 36
leukemia cutis rash cleared | 36
COVID-19 PCR became negative | 42
high-dose cytarabine consolidation | 42
tixagevimab/cilgavimab | 42
COVID-19 prophylaxis | 42
allogeneic hematopoietic stem cell transplantation | 42