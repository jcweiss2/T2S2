58 years old | 0
male | 0
hypertensive | 0
admitted to the hospital | 0
acute pancreatitis | 0
biliary or toxonutritive etiology of the pancreatitis not established | 0
WBC 12.79 | 0
BILI 19 | 0
RBC 5.31 | 0
AMS 22.38 | 0
HGB 164 | 0
AST 0.55 | 0
HCT 0.491 | 0
ALT 0.56 | 0
PLT 188 | 0
ALP 1.29 | 0
CRP 3.43 | 0
mass in the head of the pancreas 34 mm × 34 mm | 0
oncomarkers without pathological values | 0
PET-CT examination confirmed a lesion in the head of the pancreas 33 mm × 26 mm × 29 mm accumulating 16-FDG | 0
diagnosis of tumor of the pancreatic head | 0
preoperatively T2N0M0 | 0
surgical resection recommended | 0
pancreatoduodenectomy performed | 0
pancreatic duct thin | 0
pancreas had a fine structure, without fibrous component | 0
blood loss perioperatively 400 ml | 0
antibiotic prophylaxis administered | 0
octreotide administered | 0
nutrition p.o. started | 0
secretion from the drains minimal volume, without amylases | 0
drains removed on the 6th postoperative day | 0
histology findings moderately differentiated ductal adenocarcinoma pT3N0M0 with perineural invasion | 0
discharged from the hospital on the 11th postoperative day | 216
postoperative complications classified as grade II | 216
WBC 14.85 | 216
RBC 4.47 | 216
HGB 136 | 216
HCT 0.38 | 216
PLT 287 | 216
proton pump inhibitor administration started | 216
substitution of exocrine secretion of the pancreas started | 216
follow-up on the 16th postoperative day | 240
felt good, without any problems, realimented | 240
sudden upper abdominal pain appeared | 288
chills, shivers, and nausea | 288
HGB 112 | 288
RBC 3.84 | 288
WBC 10.6 | 288
HCT 0.32 | 288
PLT 483 | 288
BILI 12.7 | 288
AMS 4.25 | 288
CRP 55 | 288
ALT 0.8 | 288
AST 1.77 | 288
ALP 3.47 | 288
Q 64% | 288
INR 1.39 | 288
aPTT 24.8 | 288
spasmolytics and analgesics administered | 288
melena appeared | 288
esophagogastroduodenoscopy revealed subcardial erosions, digested blood in the stomach, coagula, and stagnation fluid | 288
acute bleeding not seen | 288
blood transfusions and i.v. antiulcer therapy administered | 288
computed tomography revealed a mass adjoining the stump of the gastroduodenal artery | 288
CT angiography of the abdominal aorta performed | 288
pseudoaneurysm of the stump of the gastroduodenal artery discovered | 288
angiography of the splanchnic arterial system confirmed bleeding from the stump of the gastroduodenal artery | 288
embolization of the gastroduodenal artery stump considered | 288
implantation of a stent graft into the common hepatic artery considered | 288
surgical procedure with resection of the bleeding pseudoaneurysm and ligation of the gastroduodenal artery stump considered | 288
implantation of a stent graft selected | 288
Jostent peripheral stent graft implanted | 288
patient under observation at the intensive care unit | 288
no signs of continued hemorrhage | 288
vital signs stable | 288
melena ceased | 288
follow-up endoscopy showed no signs of hemorrhage in the upper gastrointestinal tract | 288
antiaggregation therapy administered | 288
clopidogrel added to the patient's chronic medication | 288
7 blood transfusions administered within 48 h | 288
patient discharged | 336
postoperative radiochemotherapy completed according to plan | 720
without any problems | 720
one year after the surgery and after stent implantation | 8760