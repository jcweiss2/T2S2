40 years old | 0
man | 0
presented to the hospital | 0
hematemesis | 0
catheter ablation of the left atrium | -672
medically refractory rapid atrial fibrillation | -672
pleuritic chest pain | -504
odynophagia | -504
malaise | -504
headache | -504
fevers | -504
sepsis | 0
temperature of 100.8°F | 0
heart rate 96 bpm | 0
blood pressure 89/50 mm Hg | 0
fluid resuscitation | 0
thoracic CT with intravenous contrast | 0
small locules of gas along the esophageal wall abutting the left atrium | 0
no definite esophageal perforation | 0
no atrioesophageal fistula | 0
clinical suspicion for atrioesophageal fistula |
