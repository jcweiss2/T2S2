51 years old | 0
male | 0
admitted to the hospital | 0
moderate to severe mitral stenosis | -720
mild to moderate regurgitation | -720
atrial fibrillation | -720
chest tightness | -720
diarrhoea | -72
anti-diarrhoea medication | -72
fever | 48
high fever | 216
temperature of 38.6°C | 216
heart rate of 170 bpm | 216
blood pressure of 90/60 mmHg | 216
respiratory rate of 25 cpm | 216
slurred speech | 48
shallow left nasolabial fold | 48
grade 4 muscle strength in the left limb | 48
acute cerebral infarction | 48
cerebral haemorrhage | 48
septic shock | 216
L. adecarboxylata infection | 216
positive blood culture | 216
vegetation on the anterior leaflet of mitral valve | 216
mitral valve replacement | 240
tricuspid valvuloplasty | 240
radiofrequency ablation of atrial fibrillation | 240
left atrial auricular resection | 240
vancomycin | 216
piperacillin tazobactam | 240
levosimendan | 216
norepinephrine | 216
warfarin | 240
discharged | 720
normal biologic valve function | 720
no abnormal echogenicity around the valve | 720