26 years old | 0
man | 0
presented | 0
fever | -72
right lower limb pain | -72
swelling | -72
morbidly obese | 0
BMI 55 kg/m² | 0
gross swelling of entire right lower limb | 0
heart rate 111 beats per minute | 0
temperature 38°C | 0
leukocytosis | 0
hyperglycemia | 0
newly diagnosed type 2 diabetes mellitus | 0
source of infection not adequately removed | 0
extensive wound debridement | 0
above knee amputation | 72
ICU admission | 72
procedure uneventful | 72
required vasopressor | 72
acute renal failure | 72
metabolic acidosis | 72
swab culture obtained in OT | 72
Pseudomonas aeruginosa sensitive to amikacin | 72
gentamicin | 72
ciprofloxacin | 72
imipenem | 72
meropenem | 72
piperacillin-tazobactam | 72
cefepime | 72
imipenem-cilastatin 500 mg every 6h | 72
clindamycin 900 mg every 8h | 72
daily hemodialysis | 72
deteriorated | 72
septic shock | 72
multi-organ failure | 72
death | 120
