16 years old| 0
female | 0
fever | -336
fever (39°C, 102.2°F) | -336
generalized weakness | -336
joint pain | -336
joint pain in elbows | -336
joint pain in back | -336
auricular perichondritis | 0
ears red | 0
ears swollen | 0
joint line tenderness in elbows | 0
joint line tenderness in back | 0
joint line tenderness in multiple costochondral joints | 0
splenomegaly | 0
temperature 39°C | 0
pulse rate 102 BPM | 0
blood pressure 102/80 mmHg | 0
respiratory rate 18 respirations per minute | 0
oxygen saturation 98% | 0
hemoglobin 11.9 g/dL | 0
mean corpuscular volume 79.2 mm3 | 0
platelets 308,000/mm3 | 0
white blood cell count 14,600/mm3 | 0
CRP 369 mg/L | 0
ESR 110 mm/hr | 0
lactate dehydrogenase 561 U/L | 0
treated for suspected sepsis | 0
broad spectrum antibiotics | 0
intravenous fluids | 0
paracetamol | 0
Brucella antibodies negative | 0
cytomegalovirus negative | 0
Epstein-Barr virus negative | 0
rheumatoid factor negative | 0
ANA negative | 0
hepatitis A immunoglobulin antibodies negative | 0
bone marrow aspirate increased monocytes | 0
bone marrow normal lymphocytes | 0
bone marrow normal plasma cells | 0
Leishmania negative | 0
abdominal ultrasound spleen 15 cm | 0
abdominal ultrasound normal liver | 0
CT scan enlarged spleen | 0
CT scan mesenteric lymph node enlargement | 0
echocardiography apical hypokinesia | 0
echocardiography moderate pulmonary hypertension 50 mmHg | 0
echocardiography moderate tricuspid regurgitation | 0
echocardiography vegetation on pulmonic valve | 0
blood film microcytic hypochromic RBC | 0
blood film Rouleax formation | 0
blood film leukocytosis with segmented neutrophils | 0
blood film occasional monoblasts | 0
transferred to hematology/oncology | 0
fever persisted | 0
tachycardia 110 bpm | 0
hypotension 90/58 mmHg | 0
leukocytosis 51,000/mm3 | 0
absolute neutrophil count 36,000/mm3 | 0
hemoglobin 7.5 g/dL | 0
CRP 240 mg/L | 0
ESR 145 mm/hr | 0
broad spectrum antibiotics again | 0
urine culture negative | 0
blood culture negative | 0
transferred to ICU | 0
ferritin 3200 ng/mL | 0
fibrinogen 1.43 mg/dL | 0
total serum bilirubin 2.7 mg/dL | 0
direct serum bilirubin 1.2 mg/dL | 0
LDH 583 U/L | 0
C.ANCA negative | 0
p-ANCA negative | 0
RF negative | 0
anti-Jo negative | 0
anti-Sjögren’s-syndrome-related antigen A and B antibodies negative | 0
anti-double-stranded DNA negative | 0
anti-smith negative | 0
anti-scl-70 antibodies negative | 0
palpable purpuric lesions | 0
bullous skin lesions | 0
skin biopsy epidermal edema | 0
skin biopsy interstitial neutrophilic infiltration | 0
no evidence of vasculitis | 0
diagnosed with RP | 0
diagnosed with HLH | 0
IV fluids | 0
packed RBCs | 0
prednisolone 60 mg | 0
IVIG | 0
hydroxyurea | 0
hydroxyurea discontinued | 0
warfarin 5 mg | 0
furosemide 40 mg | 0
cyclosporine 100 mg | 0
prednisone 60 mg | 0
remission | 0
relapsed | 672
bone marrow predominance of mono-blasts | 672
bone marrow promonocytes 60% | 672
bone marrow decreased granulocytes | 672
bone marrow hypogranular cytoplasm | 672
bone marrow Pelger-Huet cells | 672
bone marrow decreased erythrocytes | 672
bone marrow decreased megakaryocytes | 672
bone marrow M:E ratio 5:1 | 672
flow cytometry FAB AML M5b | 672
AML with myelodysplasia-related changes | 672
cytarabine 160 mg | 672
allopurinol | 672
ineligible for doxuribicin | 672
AML treatment protocol incomplete | 672
Enterococcus fecium sepsis | 672
multiorgan failure | 672
died | 672
