28 years old | 0
homeless | 0
Nepalese | 0
immigrated to the United States six years previously | -52704
presented to the emergency department | 0
six months of productive cough | -4320
weight loss | -4320
intermittent abdominal pain | -4320
grade 3/6 systolic murmur heard at the right sternal border | 0
elevated hepatic transaminases | 0
computed tomography (CT) of the chest showed bilateral pleural effusions | 0
CT of the abdomen and pelvis were normal | 0
general surgery consultation obtained | 0
infectious disease consultation obtained | 0
antibiotics not given | 0
surgical intervention not recommended | 0
transthoracic echocardiogram (TTE) showed normal ejection fraction (EF) of 50–55% | 0
mobile vegetation attached to the pulmonary valve | 0
pulmonary insufficiency | 0
elevated right heart pressures | 0
bulky lesions attached to the aortic valve | 0
moderate to severe aortic insufficiency | 0
decompensated | 168
developed cardiogenic shock | 168
developed septic shock | 168
developed acute hypoxic respiratory failure | 168
treated with intravenous vancomycin | 168
treated with ceftriaxone | 168
transferred to a tertiary care facility | 168
multi-organ failure | 168
increased serum lactate level | 168
worsening oliguria | 168
initiation of continuous renal replacement therapy (CRRT) | 168
worsening clinical course | 168
hemodynamic instability | 168
high-risk surgical candidate | 168
decision to medically stabilize before surgery | 168
serology performed | 168
molecular testing performed | 168
QuantiFERON-TB Gold In-Tube testing showed latent tuberculosis infection | 168
chest x-ray not consistent with active tuberculosis | 168
three sputum specimens negative for acid-fast bacilli | 168
serology positive for Bartonella henselae IgM | 168
serology positive for Bartonella henselae IgG | 168
serology positive for Bartonella quintana IgM | 168
serology positive for Bartonella quintana IgG | 168
intravenous doxycycline treatment began on hospital day 13 | 312
gentamicin treatment began on hospital day 13 | 312
two out of 33 blood cultures positive | 2880
Candida albicans grown at two months | 1296
treated with intravenous micafungin | 1296
medical optimization for 43 days | 1032
mechanical aortic valve replacement | 1032
mitral valve repair | 1032
tissue obtained from aortic and mitral valves | 1032
16S rRNA PCR of aortic valve tissue positive for Bartonella quintana | 1032
histopathology showed vegetations | 1032
destruction of valve tissue | 1032
fibrinoid necrosis | 1032
inflammation | 1032
Warthin-Starry silver stain negative | 1032
peri-aortic thrombosis | 1032
surgical wound dehiscence | 1032
multiple thoracotomies | 1032
died | 2928
postoperative hemothorax | 2928
gastrointestinal bleeding | 2928
hemorrhagic shock | 2928
culture-negative Bartonella quintana endocarditis | 1032
history of homelessness | -52704
exposure to lice | -52704
latent tuberculosis infection | 168
no active pulmonary tuberculosis | 168
negative acid-fast bacilli on smear and culture | 168
positive QuantiFERON-TB Gold In-Tube | 168
positive respiratory syncytial virus A | 168
positive Epstein Barr virus PCR | 168
positive HSV1 PCR | 168
positive hepatitis A virus antibody (HAV Ab) | 168
positive hepatitis B surface antibody (HBsAb) | 168
negative hepatitis B surface antigen (HBsAg) | 168
negative hepatitis B core antibody (HBcAb) | 168
negative hepatitis C virus antibody (HCV Ab) | 168
cytomegalovirus PCR positive | 168
negative influenza PCR | 168
negative RMSF IgM | 168
negative Coxiella burnetti serology | 168
negative Brucella antibody | 168
negative Mycoplasma pneumonia PCR | 168
negative urine Legionella antigen | 168
