37 years old | 0
female | 0
Caucasian | 0
admitted to the hospital | 0
shortness of breath | -672
dyspnoea on exertion | -672
3rd pregnancy | -672
one healthy child | -1344
one abortion | -1344
acute toxoplasmosis | -1344
initial presentation | 0
primary care facility | 0
Bad Langensalza | 0
clinical deterioration | 0
WHO functional Class IV | 0
pulmonary embolism ruled out | 0
echocardiographic diagnosis of severe pulmonary hypertension | 0
estimated systolic PA pressure 100 mmHg | 0
transfer to intensive care unit | 0
University hospital Jena | 0
initiation of Sildenafil medication | 0
symptomatic improvement | 24
estimated systolic PA-pressure lowered to 55 mmHg | 24
emergent caesarean section | 168
stand-by mechanical circulatory support | 168
healthy child delivered | 168
transfer to standard cardiology ward | 168
right and left heart catheterization | 336
coronary artery disease ruled out | 336
arteriovenous shunts ruled out | 336
elevated mean PA pressure | 336
pulmonary vascular resistance elevated | 336
left ventricular end diastolic pressure slightly elevated | 336
secondary aetiologies ruled out | 336
diagnosis of idiopathic pulmonary hypertension | 336
sequential therapy with Macitentan initiated | 336
discharge from hospital | 720
out-patient follow-up | 1248
symptomatic patient | 1248
WHO functional Class III | 1248
elevated systolic PA pressure | 1248
right heart catheterization with vasodilator testing | 1872
elevated mean PA pressure | 1872
pulmonary vascular resistance elevated | 1872
vasodilator testing performed | 1872
significant positive result | 1872
high-dose calcium channel blocker therapy initiated | 1872
sildenafil discontinued | 1872
therapy well tolerated | 2160
symptoms improved | 2160
sequential right heart catheterization | 2160
normal values for pulmonary vascular resistance | 2160
slightly increased values for mean PA pressure | 2160
stable patient | 3024
regular out-patient visits | 3024
WHO functional class improved to I | 3024
natriuretic peptides in normal range | 3024
estimated systolic PA pressure decreased to 40 mmHg | 3024
improvements in 6 min walk test | 3024
improvements in cardiopulmonary exercise testing results | 3024
low risk | 3024
no adverse events | 3024