73 years old | 0
female | 0
arterial hypertension | -8760
calcium channel blocker | -8760
admitted to the emergency department | 0
diffuse abdominal pain | -72
right hypochondrium | -72
episodic hepatic colic | -216
fever | -168
cholestatic jaundice | -168
hemodynamically unstable | 0
blood pressure at 80/50mmgh | 0
heart rate = 135 bpm | 0
cold extremities | 0
prolonged reschooling time | 0
respiratory | 0
FR = 25 bpm | 0
SpO2 = 92% | 0
G = 1, 17 | 0
T = 39.2 | 0
BMI = 32kg/m2 | 0
oligo-anuric | 0
cardiac examination | 0
tachycardia | 0
Pleuropulmonary examination | 0
normal auscultation | 0
neurological | 0
confused | 0
GCS = 14/15th | 0
abdominal examination | 0
diffuse abdominal tenderness | 0
defense in the right hypochondrium | 0
positive murphy sign | 0
transferred to the intensive care unit | 0
conditioning | 0
vascular filling | 0
0.9% saline solution | 0
noradrenaline | 0
central venous line | 0
central venous pressure | 0
probabilistic bi-antibiotic therapy | 0
Ceftriaxon | 0
Metronidazol | 0
blood cultures | 0
electrocardiogram | 0
regular sinus rhythm | 0
HR = 137bpm | 0
transthoracic echocardiography | 0
no sign of acute cor pulmonale | 0
no disorders | 0
left ventricular ejection fraction | 0
LVEF = 50% | 0
unremarkable chest X-ray | 0
arterial blood gas | 0
uncompensated metabolic acidosis | 0
hyperlactatemia | 0
NFS | 0
leukocytosis | 0
platelet count | 0
hemoglobin | 0
inflammatory assessment | 0
CRP = 336mg/l | 0
PCT = 45 μg/l | 0
Ferritin = 1500 μg/l | 0
hemostasis assessment | 0
TP = 50% | 0
TCA | 0
hepatic assessment | 0
ASAT = 73UI/l | 0
ALAT = 92 UI/l | 0
BT = 27mg/l | 0
BD = 22mg/l | 0
GGT = 498 UI/l | 0
PAL = 425 UI/l | 0
LDH = 214UI/l | 0
urea = 4.5g/l | 0
creatinine = 100mg/l | 0
ionogram | 0
K = 7.2mEq/l | 0
Na = 137 mEq/l | 0
corrected Ca = 90mg/l | 0
lipasemia = 12 IU/l | 0
ECBU sterile | 0
abdominal ultrasound | 0
distended gallbladder | 0
thickened wall | 0
dilation of the intrahepatic bile ducts | 0
obstacle | 0
abdominal CT scan | 0
thickening of the gallbladder wall | 0
Mirizzi's SD | 0
vitamin K | 0
acute febrile Angiocholitis | 0
septic shock | 0
acute renal failure | 0
ictero-uremigenic Angiocholitis | 0
norepinephrine | 0
dobutamine | 0
hemodialysis | 24
cardiorespiratory arrest | 30
death | 30