70 years old | 0
male | 0
hypoesthesia in the fingers of each hand | -672
proximal paresis of both legs | -672
motor strength 2/5 | -672
dysfunction of gait and standing | -672
bladder incontinence | -672
rheumatoid arthritis | -672
asthma | -672
osteoporosis | -672
admitted to the hospital | 0
ventral fusion and osteosynthetic stabilization | 24
induction of anaesthesia | 24
propofol | 24
sufentanil | 24
mask ventilation | 24
rocuronium | 24
direct laryngoscopy | 24
oral intubation | 24
Cormack–Lehane grade 1 | 24
unremarkable oropharyngeal anatomy | 24
intra-operative course of general anaesthesia | 24
tracheal tube cuff pressure measurement | 24
cuff pressure briefly approached critical values | 24
spreading of tissues | 24
splitting of the sternocleidomastoid muscle compartment | 24
lateral displacement of carotid sheath | 24
microdiscectomy | 24
PEEK cage fusion | 24
osteosynthetic stabilisation | 24
unusually large hyoid bone | 24
swelling of the left side of the throat | 195
suspicion of surgery-induced hematoma | 195
laryngeal structures could be clearly palpated | 195
postponed extubation | 195
computed tomography scan | 195
cervical spine CT scan | 195
3D reconstruction | 195
fixation of the right dorsal portion of the hyoid bone | 195
fixation of the right superior horn of the thyroid cartilage | 195
leftward dislocation of the entire larynx | 195
large hematoma was ruled out | 195
transferred to the neurosurgical intensive care unit | 195
referred for Otolaryngology opinion | 195
attempt at endolaryngeal repositioning | 216
microlaryngoscopy | 216
constant readiness to perform a tracheotomy | 216
open repositioning | 240
reopening the wound | 240
hyoid bone spontaneously released | 240
CT scan | 240
normal position of the laryngeal cartilage | 240
substantial oedema | 240
mucous membranes tightly surrounded the endotracheal tube | 240
anti-oedema therapy with dexamethasone | 240
extubation | 144
respiratory insufficiency | 150
reintubation | 150
bilateral pleural effusions | 150
decreasing level of consciousness | 150
non-invasive ventilation | 150
oral reintubation | 150
unremarkable oropharyngeal anatomy | 150
conventional open tracheotomy | 288
septic | 300
ventilator-associated pneumonia | 300
antibiotic therapy | 300
reducing the level of sedation | 300
decreased level of consciousness | 300
neurological improvement was slow | 300
discharged into neurological early rehabilitation | 696
awake and oriented | 696
followed simple commands | 696
breathing using the T-piece | 696