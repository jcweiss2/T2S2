72 years old | 0
female | 0
hypothyroidism | 0
hyperlipidemia | 0
hypertension | 0
osteoarthritis | 0
severe abdominal pain | -8
vaginal bleeding | -8
bilateral oophorectomy | -960
ovarian cysts | -960
bilateral knee replacements | -960
colonoscopy | -17520
benign findings | -17520
severe nausea | 0
vomiting | 0
chills | 0
denied fever | 0
denied changes in bowel habits | 0
denied pain when urinating | 0
temperature 98.4°F | 0
blood pressure 128/84 mmHg | 0
heart rate 104 bpm | 0
respiration rate 20 breaths per minute | 0
O2 saturation 98% | 0
severe distress | 0
tympanic distended abdomen | 0
tender to palpation | 0
rebound tenderness | 0
moderate leukocytosis (12600/mm3) | 0
anion gap metabolic acidosis | 0
bicarbonate 15 | 0
azotemia | 0
BUN 26 | 0
creatinine 2.6 mg/dL |7 0
Foley catheter placement | 0
minimal urine output | 0
2 L normal saline administration | 0
gynecology consultation | 0
uterine prolapse | 0
mild vaginal bleeding | 0
CT abdomen and pelvis with contrast | 0
pneumoperitoneum | 0
pneumobilia | 0
large masslike collection of mottled air and soft-tissue density | 0
suggesting intrauterine infection or necrosis | 0
colonic perforation | 0
possible enterofistula connecting to the uterus | 0
no evidence of obstruction | 0
no other signs of inflammatory disease | 0
exploratory laparotomy | 0
foul-smelling gas burst | 0
2.5 cm spontaneous rupture of posterior fundus | 0
suspected intrauterine malignancy | 0
total abdominal hysterectomy | 0
salpingectomy | 0
mass on distal appendix | 0
appendectomy | 0
small bowel examination | 0
colon examination | 0
peritoneal cavity irrigation with normal saline | 0
antibiotic solution irrigation | 0
peritoneal-cavity fluid cultures | 0
uterine myometrial tissue pathology | 0
abdomen closure with retention sutures | 0
Jackson-Pratt drain placement | 0
severe end organ damage | 0
multi end organ failure | 0
intubated | 0
transfer to surgical ICU | 0
advanced high-grade serous adenocarcinoma of the endometrium | 0
>50% invasion into myometrium | 0
blood gram stain showing gram-positive rods | 0
C. perfringens confirmed by blood cultures | 0
intraoperative wound cultures | 0
POD 0 | 0
severely acidemic | 0
hypotensive | 0
norepinephrine administration | 0
broad-spectrum antibiotics (piperacillin/tazobactam, vancomycin, metronidazole) | 0
POD 1 | 24
positive C. perfringens in blood and peritoneal fluid cultures | 24
antibiotic regimen changed to vancomycin and IV penicillin G | 24
POD 4 | 96
abdomen increasingly tense and distended | 96
worsening multiorgan failure secondary to sepsis | 96
reexploration of abdominal cavity | 96
large quantity of brown and ashy fluid removed | 96
necrosis of distal half of small bowel | 96
necrosis of entire colon | 96
necrosis of proximal rectum | 96
ileectomy | 96
total colectomy | 96
proximal rectum resection | 96
peritoneal cavity washout | 96
bowel left in discontinuity | 96
wound vacuum placement | 96
POD 6 | 144
ileostomy creation | 144
focal areas of patchy necrosis at 5 small bowel sites | 144
contiguous resection not possible | 144
multiple resections | 144
ileostomy created | 144
postoperative necrosis at ileostomy site | 144
hemodynamic instability | 144
advance directives revisited with family | 144
comfort care with terminal wean | 144
patient died | 144
