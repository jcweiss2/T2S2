32 years old | 0
Gravida 2 Para 2 | 0
admitted to the hospital | 0
fevers | -168
chills | -168
left distal lower extremity pain | -168
left distal lower extremity swelling | -168
right knee swelling | -168
diffuse rash | -168
denies recent injury | -168
unable to bear weight on the left side | -168
continued breastfeeding | -168
history of stage IIa malignant peripheral nerve sheath tumor | -8760
treated 1-year prior | -8760
complete surgical excision | -8760
no chemotherapy | -8760
admitted in labor | -168
420/7 weeks gestation | -168
uncomplicated antepartum course | -168
group B streptococcus carrier screening negative | -168
small labial and first-degree midline lacerations | -168
repaired at time of delivery | -168
minimal blood loss | -168
discharged home on postpartum day 1 | -144
fevers to 104°F at home | -144
temperature 97.5°F | 0
heart rate 68 bpm | 0
respiratory rate 18 | 0
blood pressure 107/69 | 0
mild distress | 0
moderate pain | 0
limited range of motion of the left lower extremity | 0
focal area of erythema | 0
exquisitely tender to palpation | 0
right knee swollen | 0
peripheral pulses present | 0
abdomen nonperitoneal | 0
uterus mildly tender | 0
fundus firm at 4-cm below the umbilicus | 0
faint maculopapular rash | 0
scant nonpurulent lochia | 0
leukocytosis to 18,800 | 0
bandemia of 23.7% | 0
lactate of 1.6% | 0
clean-catch urine culture positive for S. pyogenesis | 0
orthopaedics consulted | 0
concern for possible compartment syndrome | 0
concern for underlying GAS necrotizing infection | 0
plain X-ray films demonstrated soft tissue edema | 2
Doppler ultrasonography negative for deep vein thrombosis | 2
left ankle arthrocentesis performed | 2
normal appearing fluid obtained | 2
vital signs notable for HR = 144 bpm | 2
T = 102.6°F | 2
RR = 20 | 2
MAP = 66 | 2
SpO2 = 98% | 2
aggressive fluid resuscitation initiated | 2
blood cultures obtained | 2
IV amoxicillin-sulbactam and clindamycin started | 2
transfer to ICU | 2
CT of the left lower extremity noted severe inflammation | 4
left distal lower extremity anterior and lateral compartment fasciotomy | 6
no purulence or necrotic tissue noted | 6
normal appearing fascia | 6
improvement in pain | 6
albumin administered | 6
norepinephrine administered | 6
esmolol administered | 6
gentamicin administered | 6
therapeutic enoxaparin administered | 6
tachycardia resolved | 120
fevers resolved | 120
leukocytosis resolved | 120
stable for transfer out of ICU | 120
residual peroneal nerve palsy | 192
reoperation of the left distal lower extremity | 192
concerns of myositis | 192
small area of purulence | 192
decreased contractility of the anterior compartment | 192
fever to 102.2°F | 312
new leukocytosis | 312
worsening pain in right knee | 312
arthrocentesis performed | 312
frank purulent fluid obtained | 312
right knee arthroscopy | 312
synovectomy and debridement | 312
inflamed proliferative synovium | 312
repeat right knee arthroscopic incision and drainage | 336
negative culture | 336
transitioned to IV penicillin G | 408
discharged to home | 456
continued treatment with IV penicillin | 456
follow-up visits with orthopaedics | 480
no evidence of osteomyelitis | 480
no continued infection | 480
chondromalacia of left patella diagnosed | 480
persistent residual peroneal palsy | 480
poor wound healing | 480
multiple enlarged inguinal lymph nodes | 480
enlargement on ultrasound | 504
reactive process suspected | 504
left inguinal lymph node excisional biopsy | 744
left lower leg wound debridement | 744
lymph node biopsy negative for metastatic tumor | 744
reactive follicular hyperplasia | 744
final blood cultures and infectious laboratories confirmed resolution of GAS infection | 744