32 years old | 0
female | 0
intravenous drug use | -672
attention deficit/hyperactivity disorder | -672
fever | -168
chills | -168
generalized weakness | -168
shortness of breath | -72
admitted to the hospital | 0
temperature 102.7 °Fahrenheit | 0
blood pressure 102/56 mmHg | 0
pulse 136 beats per minute | 0
respiratory rate 38 breaths per minute | 0
oxygen saturation 94% | 0
bilateral rhonchi | 0
tachycardia | 0
no murmur | 0
no rub | 0
no gallop | 0
WBC 12,200/mm3 | 0
hemoglobin 10.9 g/dL | 0
platelet count 85,000/mm3 | 0
ESR 60 mm/hr | 0
hyponatremia | 0
sodium 124 mmol/L | 0
creatinine level 2.8 mg/dL | 0
BUN 98 mg/dL | 0
NT-proBNP 1028 pg/mL | 0
sinus tachycardia | 0
bilateral lower lobe infiltrates | 0
small pleural effusions | 0
given IV fluids | 0
given levofloxacin | 0
clinical condition deteriorated | 24
transferred to ICU | 24
septic shock | 24
acute respiratory failure | 24
pressor support | 24
mechanical ventilation | 24
blood cultures grew gram-positive cocci | 24
started vancomycin | 24
tricuspid valve vegetation | 48
moderate-to-severe tricuspid regurgitation | 48
patent foramen ovale | 48
shunt | 48
multiple cavitary peripheral lung nodules | 48
septic emboli | 48
non-oliguric AKI | 48
renal replacement therapy | 48
acute tubular necrosis | 48
MSSA | 72
started oxacillin | 72
improved on supportive and antimicrobial therapy | 168
weaned off pressors | 168
extubated | 168
renal function recovered | 168
skin examination revealed bilateral nontender purpuric papules | 216
palpable purpuric papules | 216
bullous lesions | 240
no mucosal involvement | 216
no palmar involvement | 216
no abdominal pain | 216
no arthralgias | 216
no paresthesia | 216
no fever | 216
no chills | 216
HIV antibody negative | 216
hepatitis B serology negative | 216
p-ANCA negative | 216
c-ANCA negative | 216
cryoglobulin negative | 216
rheumatoid factor negative | 216
ANA weakly positive | 216
anti-ds DNA antibody negative | 216
complement C3 low | 216
complement C4 normal | 216
anti-HCV antibody positive | 216
HCV viral load 4.16 × 105 IU/mL | 216
eosinophil count normal | 216
aspirated fluid from bullous lesions did not grow bacteria | 240
no organisms seen on gram staining | 240
punch biopsies from bullous skin lesions showed perivascular neutrophil infiltration | 240
fibrinoid necrosis of small vessels | 240
leukocytoclastic vasculitis | 240
vancomycin started | 240
oxacillin discontinued | 240
skin lesions resolved | 312
tricuspid valve replacement surgery | 720
no perioperative complications | 720
follow-up appointment | 720
no recurrence of skin lesions | 720