63 years old | 0
    woman | 0
    acute onset fever | 0
    chills | 0
    malaise | 0
    cigarette smoking | 0
    previous breast cancer resection | 0
    dog hand bite | -48
    creatinine 1.22 mg/dl | 0
    lactate dehydrogenase 298 | 0
    AST 115 | 0
    ALT 54 U/l | 0
    hyponatremia 130 mmol/l | 0
    hyposmolality 265 mOsm/kg | 0
    PaO2/FiO2 ratio 246 mmHg | 0
    bilateral basal hyperdensities of the lungs | 0
    admitted to the medicine department | 0
    diagnosis of pneumonia | 0
    empirical antibiotic therapy with levofloxacin | 0
    thrombocytopenia | 24
    acute kidney injury | 24
    livedo reticularis | 24
    arterial hypotension | 24
    acute hypoxemic respiratory failure | 24
    high serum procalcitonin 79.7 ng/ml | 24
    Gram-negative rods in blood culture | 24
    empirical course of meropenem | 24
    admitted to the ICU | 24
    intubated | 24
    condition worsened to full-blown septic shock | 24
    severe lactic acidosis | 24
    high-dose inotropic support | 24
    continuous mandatory mechanical ventilation | 24
    hydrocortisone 200 mg/die | 24
    AKI stage 3 | 24
    anuria | 24
    serum creatinine 3.91 mg/dl | 24
    renal replacement therapy | 24
    rhabdomyolysis | 96
    liver injury | 96
    severe thrombocytopenia | 96
    coagulopathy | 96
    fresh frozen plasma transfusion | 96
    platelet transfusion | 96
    livedo reticularis worsened to frank purpura | 96
    ischemia of the limbs | 96
    blood culture became positive | 168
    microbiological diagnosis of C. canimorsus | 168
    started ampicillin-sulbactam | 168
    started ceftriaxone | 168
    resolution of critical illness | 168
    isolated strain sensitive to multiple antibiotics | 168
    surgical amputation of finger | 336
    surgical amputation of inferior limbs below knees | 336
    end-stage renal disease | 336
    intermittent hemodialysis | 336
    