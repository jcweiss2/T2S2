32 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
intravenous drug use | -672 | 0 | Factual
attention deficit/hyperactivity disorder | -672 | 0 | Factual
fevers | -168 | 0 | Factual
chills | -168 | 0 | Factual
generalized weakness | -168 | 0 | Factual
shortness of breath | -72 | 0 | Factual
abusing fentanyl intravenously | -672 | 0 | Factual
dextroamphetamine/amphetamine | -672 | 0 | Factual
no exposure to other medications or chemicals | 0 | 0 | Factual
admitted to the hospital | 0 | 0 | Factual
Temperature 102.7 °Fahrenheit | 0 | 0 | Factual
blood pressure 102/56 mmHg | 0 | 0 | Factual
pulse 136 beats per minute | 0 | 0 | Factual
respiratory rate 38 breaths per minute | 0 | 0 | Factual
oxygen saturation 94% on room air | 0 | 0 | Factual
moderate respiratory distress | 0 | 0 | Factual
bilateral rhonchi | 0 | 0 | Factual
tachycardia | 0 | 0 | Factual
no murmur, rub or gallop | 0 | 0 | Negated
WBC 12,200/mm3 | 0 | 0 | Factual
hemoglobin 10.9 g/dL | 0 | 0 | Factual
platelet count 85,000/mm3 | 0 | 0 | Factual
ESR 60 mm/hr | 0 | 0 | Factual
hyponatremia with sodium 124 mmol/L | 0 | 0 | Factual
creatinine level 2.8 mg/dL | 0 | 0 | Factual
BUN 98 mg/dL | 0 | 0 | Factual
NT-proBNP 1028 pg/mL | 0 | 0 | Factual
sinus tachycardia | 0 | 0 | Factual
bilateral lower lobe infiltrates | 0 | 0 | Factual
small pleural effusions | 0 | 0 | Factual
given IV fluids | 0 | 24 | Factual
levofloxacin intravenously | 0 | 24 | Factual
septic shock | 24 | 24 | Factual
acute respiratory failure | 24 | 24 | Factual
pressor support | 24 | 168 | Factual
mechanical ventilation | 24 | 168 | Factual
blood cultures grew gram-positive cocci | 24 | 24 | Factual
vancomycin therapy | 24 | 168 | Factual
tricuspid valve vegetation | 48 | 48 | Factual
moderate-to-severe tricuspid regurgitation | 48 | 48 | Factual
patent foramen ovale with shunt | 48 | 48 | Factual
septic emboli | 48 | 48 | Factual
non-oliguric AKI | 48 | 168 | Factual
renal replacement therapy | 48 | 168 | Factual
MSSA | 72 | 72 | Factual
oxacillin treatment | 72 | 240 | Factual
improved on supportive and antimicrobial therapy | 168 | 240 | Factual
weaned off pressors | 168 | 240 | Factual
extubated | 168 | 240 | Factual
renal function recovered | 168 | 240 | Factual
skin examination revealed bilateral nontender purpuric papules | 240 | 240 | Factual
bullous lesions | 264 | 288 | Factual
no mucosal or palmar involvement | 240 | 288 | Negated
no abdominal pain | 240 | 288 | Negated
no arthralgias | 240 | 288 | Negated
no paresthesia | 240 | 288 | Negated
no fever | 240 | 288 | Negated
no chills | 240 | 288 | Negated
HIV antibody negative | 240 | 240 | Factual
hepatitis B serology negative | 240 | 240 | Factual
p-ANCA negative | 240 | 240 | Factual
c-ANCA negative | 240 | 240 | Factual
cryoglobulin negative | 240 | 240 | Factual
rheumatoid factor negative | 240 | 240 | Factual
ANA weakly positive | 240 | 240 | Factual
anti-ds DNA antibody negative | 240 | 240 | Factual
Complement C3 low | 240 | 240 | Factual
Complement C4 normal | 240 | 240 | Factual
anti-HCV antibody positive | 240 | 240 | Factual
HCV viral load 4.16 × 105 IU/mL | 240 | 240 | Factual
eosinophil count normal | 240 | 288 | Factual
aspirated fluid from bullous lesions did not grow bacteria | 264 | 264 | Factual
no organisms seen on gram staining | 264 | 264 | Factual
punch biopsies from bullous skin lesions showed perivascular neutrophil infiltration | 264 | 264 | Factual
fibrinoid necrosis of small vessels | 264 | 264 | Factual
leukocytoclastic vasculitis | 264 | 264 | Factual
vancomycin started in lieu of oxacillin | 288 | 288 | Factual
resolution of skin lesions | 288 | 720 | Factual
tricuspid valve replacement surgery | 720 | 720 | Factual
no recurrence of skin lesions | 720 | 720 | Factual