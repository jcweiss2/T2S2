seven years old | 0 | 0 
male | 0 | 0 
admitted to the hospital | 0 | 0 
pre-B-ALL | -672 | 0 
first relapse of pre-B-ALL | -336 | -168 
allogeneic HSCT | -168 | -168 
second relapse of pre-B-ALL | -24 | 0 
hemoglobin 8.5 g/dl | 0 | 0 
thrombocytes 13,000/μl | 0 | 0 
WBC 940/μl | 0 | 0 
neutrophils 50/μl | 0 | 0 
CRP 6.83 mg/dl | 0 | 0 
ferritin 182 μg/dl | 0 | 0 
cachexia | 0 | 0 
dry skin | 0 | 0 
pallor | 0 | 0 
multiple hematomas | 0 | 0 
hepatosplenomegaly | 0 | 0 
antibiotic, antiviral, and antifungal chemoprophylaxis | 0 | 168 
ceftriaxone | 0 | 168 
teicoplanin | 0 | 168 
acyclovir | 0 | 168 
caspofungin | 0 | 168 
pain in the left flank | -24 | 0 
morphine | -24 | 120 
blinatumomab treatment | 0 | 168 
aggravation of pain | 120 | 120 
somnolent and sleepy | 144 | 144 
cerebral side effect of blinatumomab | 144 | 144 
neurological condition worsened | 144 | 168 
cerebral CT scan | 144 | 144 
MRI scan | 144 | 144 
multiple cerebral hemorrhages | 144 | 168 
cardio-respiratory decompensation | 168 | 168 
mechanical ventilation | 168 | 168 
catecholamine therapy | 168 | 168 
blinatumomab treatment stopped | 168 | 168 
hemoglobin 6.7 g/dl | 168 | 168 
thrombocytes 49,000/μl | 168 | 168 
WBC 120/μl | 168 | 168 
neutrophils 20/μl | 168 | 168 
CRP 23.13 mg/dl | 168 | 168 
ferritin 1439 μg/dl | 168 | 168 
multiple thrombi in the left and right ventricle | 168 | 168 
thromboembolic events | 168 | 168 
endocarditis | 168 | 168 
septic embolisms | 168 | 168 
meropenem | 168 | 168 
gentamicin | 168 | 168 
CT scans of the thorax, abdomen and pelvis | 168 | 168 
multiple, systemic thromboembolic lesions | 168 | 168 
ischemia | 168 | 168 
bleeding | 168 | 168 
infarction | 168 | 168 
bone marrow aplasia | 168 | 168 
lymphatic blasts | 168 | 168 
cerebral pressure rising | 168 | 168 
cerebral herniation | 168 | 168 
death | 168 | 168 
invasive mycosis of R. pusillus | 0 | 168 
autopsy | 168 | 168 
R. pusillus identified via PCR-based methods | 168 | 168 
disseminated mucormycosis | 0 | 168 
mucormycosis in lungs | 0 | 168 
mucormycosis in other organs | 0 | 168 
health care-related infection | 0 | 168 
liposomal amphotericin B | 168 | 168 
posaconazole | 168 | 168 
breakthrough filamentous fungal infections | 168 | 168 
resistant fungi | 168 | 168 
fulminant mucormycosis during blinatumomab treatment | 0 | 168 
targeted therapy | 0 | 168 
reduced immunocompetence after HSCT | 0 | 168 
invasive fungal infections | 0 | 168 
antifungal prophylaxis | 0 | 168 
prophylactic treatment with an antimycotic medication | 168 | 168 
covering mucormycetes | 168 | 168