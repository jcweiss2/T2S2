77 years old | 0
lady | 0
ASA III | 0
scheduled for emergency laparotomy | 0
hollow viscous perforation | 0
abdominal pain | -24
fever | -24
febrile | 0
pulse 110/min | 0
regular pulse | 0
blood pressure 106/72 mmHg | 0
respiratory rate 20/min | 0
no abnormal heart sounds | 0
no abnormal breath sounds | 0
haemoglobin 11.9 g/dl | -6
total counts 14,000/mm3 | -6
band forms 13% | -6
serum sodium 140 mEq/l | -6
potassium 3.6 mEq/l | -6
platelets 220,000/mm3 | -6
creatinine 1.4 mg% | -6
bilateral mild pleural effusion | -6
sinus tachycardia | -6
heart rate 106/min | -6
ECG showed HR 156/min in AF | 0
invasive blood pressure 106/72 mmHg | 0
SpO2 93% on 60% oxygen | 0
intravenous metoprolol administered | 0
no change in HR | 0
defibrillator kept available | 0
trachea intubated | 0
rapid sequence induction | 0
midazolam 1 mg administered | 0
fentanyl 250 mcg administered | 0
propofol 60 mg administered | 0
succinylcholine 60 mg administered | 0
central line inserted | 0
anaesthesia maintained | 0
air | 0
oxygen | 0
sevoflurane | 0
fentanyl | 0
hydromorphone | 0
rocuronium | 0
intravenous amiodarone 150 mg administered | 0
HR reduced to 80-90/min | 15
improvement in blood pressure | 15
rhythm reverted back to sinus | 15
uncompensated metabolic acidosis | 15
bicarbonate 16 mEq/l | 15
respiratory alkalosis | 15
PCO2 26 mmHg | 15
serum potassium 3 mEq/l | 15
intravenous potassium 20 mmol/L administered | 15
repeat serum potassium 3.4 mEq/l | 60
intraoperative period uneventful | 120
transferred to ICU | 120
IV potassium supplementation | 120
IV magnesium sulphate administered | 120
serum magnesium 1.2 mg/dl | 120
calcium chloride administered | 120
serum calcium 6 mg/dl | 120
elevated CRP | 120
elevated procalcitonin | 120
thyroid function tests normal | 120
trachea extubated | 12
controlled ventricular rate | 12
sinus rhythm | 12
tab. aspirin 81 mg once daily started | 12
negative transthoracic echocardiogram | 12
discharged home | 168
low-dose aspirin therapy | 168