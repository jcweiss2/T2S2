77 years old | 0
male | 0
admitted to the hospital | 0
left iliac fossa pain | -72
diarrhoea | -72
nausea | -72
vomiting | -72
fevers | -72
past history of advanced prostate cancer | -6720
bony metastasis | -6720
previous chemotherapy | -6720
radiotherapy | -6720
type two diabetes mellitus | -6720
abiraterone | -6720
prednisolone | -6720
flutamide | -6720
oxycodone | -6720
targin | -6720
sinus tachycardia | 0
elevated temperature | 0
diffuse tenderness | 0
positive bowel sounds | 0
low haemoglobin | 0
low white cell count | 0
normal coagulation | 0
normal liver function | 0
normal lipase | 0
normal lactate | 0
grossly thickened small bowel | 0
portal venous gas in liver | 0
conservative treatment | 0
fluid resuscitation | 0
intravenous tazocin | 0
granulocyte-colony stimulating factor | 0
nasogastric decompression | 0
rising C-reactive protein | 24
exploratory laparotomy | 24
moderate bowel oedema | 24
no bowel or mesenteric necrosis | 24
division of adhesions of the jejunum and ileum | 24
diagnosis of chemotherapy/radiotherapy-related severe enterocolitis | 24
small bowel obstruction | 120
transferred back to the rural hospital | 648