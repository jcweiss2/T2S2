40 years old | 0
male | 0
admitted to the hospital | 0
odynophagia | -168
dry cough | -168
exertional dyspnea | -168
fever | -168
arthralgias | -168
fatigue | -168
diabetes | -6720
glycosylated hemoglobin 10.8 % | -6720
insulin treatment | -6720
glargine | -6720
lispro | -6720
body mass index 28.3 kg / m2 | 0
heart rate 110 beats per minute | 0
24 breaths per minute | 0
oxygen saturation of 82 % | 0
right lung rales | 0
no cyanosis | 0
no lower limb edema | 0
no history of smoking | 0
no alcohol consumption | 0
arterial gases showed moderate oxygen impairment | 0
supplemental oxygen required | 0
normal blood count | 0
increased CRP | 0
right basal ground glass opacity | 0
positive RT-PCR COVID- 19 | 0
adenovirus isolated | 0
lactate dehydrogenase increased | 0
ferritin markedly elevated | 0
D-dimer positive | 0
ground-glass opacities with multilobar involvement | 0
transferred to intensive care unit | 144
dyspnea increased | 144
tachypnea | 144
desaturation | 144
ampicillin-sulbactam started | 144
clarithromycin started | 144
hydroxychloroquine started | 144
hypotension developed | 144
hypoxemia developed | 144
mechanical ventilation started | 144
norepinephrine started | 144
septic shock diagnosed | 144
acute respiratory distress syndrome diagnosed | 144
pronation | 144
neuromuscular relaxation cycles | 144
Klebsiella oxytoca isolated | 144
antibiotic escalation to cefepime | 144
extubation | 432
transferred to general floor | 432
symptoms resolved | 432
second RT-PCR SARS Cov2 negative | 480
discharged | 480
supplemental oxygen requirement at home | 480