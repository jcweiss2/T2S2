35 years old | 0
male | 0
autosomal dominant polycystic kidney disease | 0
admitted to the hospital | 0
kidney transplantation | 0
methylprednisolone | 0
basiliximab | 0
rabbit anti-human thymocyte immunoglobulin (ATG) | 0
tacrolimus | 0
mycophenolate mofetil | 0
prednisone | 0
Corynebacterium detected in donor kidney preservation solution | -96
no evidence of Corynebacterium-related infection | -96
discharged | 336
low fever | 1344
light hematuria | 1344
mild frequent urination | 1344
urgent urination | 1344
painful urination | 1344
white blood cell count of 17.46×10^9/L | 1344
hemoglobin level of 95 g/L | 1344
C-reactive protein level of 231.06 mg/L | 1344
serum creatinine (Scr) level of 196.1 µmol/L | 1344
prothrombin time of 15.40 s | 1344
blood pressure of 87/64 mmHg | 1344
partial intracapsular hemorrhage in primary bilateral polycystic kidneys | 1344
septic shock | 1344
disseminated intravascular coagulation | 1344
readmitted to hospital | 1344
supportive treatment | 1344
maintenance immunosuppressive regimen tapered | 1344
mycophenolate withdrawn | 1344
tacrolimus replaced by cyclosporin | 1344
meropenem administered | 1344
Corynebacterium found in patient's blood | 1392
Enterococcus faecium found in patient's urine | 1392
Pseudomonas putida found in patient's urine | 1392
linezolid administered | 1392
ultrasound examination | 1512
no special finding | 1512
cyclosporin replaced by tacrolimus | 1512
troponin T and atrial natriuretic peptide levels increased | 1536
chest pain | 1536
dyspnea | 1536
inability to lie in supine position | 1536
electrocardiogram revealed sinus tachycardia with premature ventricular beats | 1536
acute anuria | 1536
gradual increase in Scr to 346 µmol/l | 1536
multiple thromboses found in right external iliac artery | 1536
transferred to intensive care unit | 1536
bedside continuous renal replacement therapy | 1536
adjusted scheme of meropenem and vancomycin | 1536
sudden persistent angina pectoris | 1560
chest tightness | 1560
no sweating | 1560
increase in myocardial enzymes | 1560
cardiac murmur | 1560
echocardiography revealed medium echoic mass at posterior mitral valve tip | 1560
moderate-to-severe mitral regurgitation | 1560
mild-to-moderate tricuspid regurgitation | 1560
non-ST segment elevation myocardial infarction diagnosed | 1560
fraxiparin administered | 1560
cough with bloody sputum | 1656
fraxiparin stopped | 1656
operation scheduled | 1692
allograft nephrectomy planned | 1692
mitral valve replacement and vegetative resection planned | 1692
cardiac arrest | 1692
ventricular fibrillation | 1692
emergency external chest compression | 1692
electric defibrillation | 1692
endotracheal intubation | 1692
mitral valve replacement surgery and vegetative resection performed | 1692
allograft nephrectomy not performed | 1692
large polypoid vegetation found attached to posterior leaflet of mitral valve | 1692
patient died | 1752
metagenomic next-generation sequencing (mNGS) performed | 8760
Corynebacterium striatum identified | 8760