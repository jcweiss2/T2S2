53 years old| 0
male| 0
admitted to the hospital| 0
hydronephrosis| 0
urolithiasis| 0
ureteral stent placement (left side)| 0
hypertension| -72
hypercholesterolemia| -72
violent pain in epigastric region| 72
nausea| 72
pale| 72
sweaty| 72
cold| 72
sinus tachycardia (120 beats/min)| 72
hypotension (90/70 mm Hg)| 72
distended abdomen| 72
moderate tenderness in epigastrium| 72
moderate tenderness in left hypochondrium| 72
anemia| 72
thrombopenia| 72
slight increase in international normalized ratio| 72
slight increase in activated partial thromboplastin time| 72
slight increase in alanine aminotransferase| 72
decompensated metabolic acidosis| 72
rapid resuscitation with intravenous crystalloid solutions| 72
stabilization of hemodynamic status| 72
focussed assessment with sonography for trauma scan| 72
free fluid in all recesses of peritoneal cavity| 72
contrast-enhanced CT scan of abdomen and pelvis| 72
dilated left hepatic artery| 72
bleeding point (aneurysm 20 x 18 mm)| 72
aneurysm originating from left gastric artery| 72
large intraperitoneal effusion| 72
heterogeneous hepatic enhancement in left lateral liver segments| 72
hepatic hypoperfusion| 72
laparotomy| 72
massive hemoperitoneum (1500 mL)| 72
ruptured aneurysm of hepatic arterial branch| 72
fresh blood clot in artery| 72
diffused disruption of vascular wall| 72
clamped aneurysm| 72
isolated proximal stump up to origin of left hepatic artery| 72
no clinical sign of hepatic ischemia after cross-clamping| 72
complete aneurysmectomy| 72
intensive care unit admission (first 48 hours)| 72
correction of acidosis during surgery| 72
stabilization of hemodynamic conditions| 72
transfer to surgical ward| 120
noninfectious fever| 120
hospital stay prolonged| 120
discharged from hospital| 360
asymptomatic at discharge| 360
liver function tests within normal ranges| 360
rupture of hepatic artery aneurysm| 72
hemoperitoneum| 72
replaced left hepatic artery from left gastric artery| 72
replaced right hepatic artery from superior mesenteric artery| 72
atherosclerosis (etiology)| 72
hypertension (risk factor)| 72
hypercholesterolemia (risk factor)| 72
hepatic ischemia not observed| 72
postoperative acidosis correction| 72
hemodynamic stabilization| 72
noninfectious fever onset| 120
postoperative complications| 120
discharge after 15 days| 360
