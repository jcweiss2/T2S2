72 years old | 0
male | 0
clinically quiescent Crohn's disease | -672
fever | -96
fatigue | -96
altered mental status | -96
nausea/vomiting | -96
diagnosis of acute myelogenous leukemia (AML) | -96
tumor lysis syndrome | -96
acute kidney injury (AKI) | -96
hyperleukocytosis | -96
ICU admission | -96
treated empirically with ceftazidime | -96
treated empirically with vancomycin | -96
blood cultures were sterile | -96
urine cultures were sterile | -96
CT of the chest, abdomen, and pelvis was unremarkable | -96
neutropenic | -48
cytoreductive therapy with hydroxyurea | -48
cytoreductive therapy with cytarabine | -48
dose-reduced G-CLAM | -48
defervesced | -48
ceftazidime continued | 0
vancomycin stopped | 0
fever | 0
mild abdominal pain | 24
new diarrhea | 24
enteric pathogen panel obtained | 24
Biofire FilmArray GI panel | 24
blood agar plate | 24
loperamide started | 48
MRSA detected on blood agar plate | 72
oral vancomycin started | 72
piperacillin-tazobactam started | 72
respiratory distress | 96
intubated | 96
recurrence of AKI | 96
recurrence of shock | 96
vancomycin IV added | 96
CT of the abdomen and pelvis showed diffuse small bowel wall edema | 96
CT of the abdomen and pelvis showed thickening | 96
CT of the abdomen and pelvis showed dilatation | 96
CT of the abdomen and pelvis showed pneumatosis | 96
transitioned to comfort care | 96
expired | 96
postmortem evaluation revealed gross dilatation of the duodenum and jejunum | 96
postmortem evaluation revealed dusky discoloration | 96
postmortem evaluation revealed mucosal erythema and congestion | 96
postmortem evaluation revealed Gram positive cocci | 96
focal mucosal erosions in the stomach | 96
focal mucosal erosions in the cecum | 96
no pseudomembranes found | 96
cause of death was septic shock with multiorgan failure | 96
cause of death was secondary to MRSA enterocolitis | 96