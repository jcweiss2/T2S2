73 years old | 0
male | 0
unconscious | 0
found at home | 0
brought to the emergency department by ambulance | 0
empty bottle of Supracide insecticide | 0
methidathion | 0
suicide note found | 0
past medical history unremarkable | 0
no hypertension | 0
no diabetes | 0
body weight approximately 45 kg | 0
comatose | 0
Glasgow coma scale score of 3 | 0
pupils pinpoints | 0
blood pressure 120/100 mm Hg | 0
pulse rate 108 per minute | 0
respiration rate 24 per minute | 0
body temperature 36°C | 0
salivation increased | 0
rales increased in both lung fields | 0
intubated | 0
mechanical ventilation | 0
activated charcoal given via nasogastric tube | 0
repeated boluses of atropine given in 2-mg aliquots | 0
clear lung sounds heard | 0
continuous infusion of atropine started at 1 mg/hr | 0
infusion titrated until clear breathing sounds heard | 0
infusion of pralidoxime started at 500 mg/hr | 0
arterial pH 7.220 | 0
partial pressure of carbon dioxide (PCO2) 36.7 mm Hg | 0
PO2 59.9 mm Hg | 0
bicarbonate 14.7 mmol/L | 0
serum lactate 7.8 mmol/L | 0
blood urea nitrogen 18 mg/dl | 0
serum creatinine 1.2 mg/dl | 0
plasma cholinesterase level <200 units/L | 0
blood pressure dropped to 70/40 mm Hg | -6
norepinephrine infusion started | -6
norepinephrine titrated to blood pressure | -6
urine output decreased to 25 ml/hr | -6
blood gas analysis revealed pH 7.154 | -6
PCO2 20.8 mm Hg | -6
PO2 323 mm Hg | -6
bicarbonate 7.1 mmol/L | -6
serum creatinine 1.46 mg/dl | -6
CRRT initiated | -6
oliguria | -6
acidosis | -6
unstable hemodynamic condition | -6
CRRT prescription: continuous venovenous hemodiafiltration (CVVHDF) via jugular venous catheter | -6
blood flow 120 ml/min | -6
dialysate flow 500 ml/hr | -6
substitute flow 1,000 ml/hr | -6
fluid removal 200 ml/hr | -6
total effluent flow rate 37.7 ml/kg/hr | -6
norepinephrine requirement decreased | -6
norepinephrine requirement remained between 0.09–0.13 µg/kg/min for 20 hours after CRRT initiation | -6
condition progressively deteriorated | 72
maximal ventilatory support | 72
maximal hemodynamic support | 72
maximal renal support | 72
antidote therapy | 72
died | 96
plasma cholinesterase levels measured on second and third days | 24
prefilter plasma cholinesterase levels <200 U/L | 24
postfilter plasma cholinesterase 358 U/L 1 hour after CRRT initiation | -5
postfilter plasma cholinesterase 689 U/L 18 hours after CRRT initiation | 12
