42 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
admitted to the hospital | 0 | 0 | Factual
altered mental status | 0 | 0 | Factual
low grade fevers | -120 | 0 | Factual
sudden deterioration in mental status | 0 | 0 | Factual
history of intravenous drug use | -8760 | -720 | Factual
extraction of all maxillary teeth | -2160 | -2160 | Factual
mandibular dental infection | -1296 | -1296 | Factual
treated with oral amoxicillin | -1296 | -1296 | Factual
temperature was 36.7 °C | 0 | 0 | Factual
heart rate was 98 beats/min | 0 | 0 | Factual
respiratory rate was 17 breaths/min | 0 | 0 | Factual
blood pressure was 131/66 mm Hg | 0 | 0 | Factual
oxygen saturation of 99% on room air | 0 | 0 | Factual
denies fevers | 0 | 0 | Negated
denies chills | 0 | 0 | Negated
denies chest pain | 0 | 0 | Negated
denies dyspnea | 0 | 0 | Negated
denies nausea | 0 | 0 | Negated
denies vomiting | 0 | 0 | Negated
denies diarrhea | 0 | 0 | Negated
denies skin lesions | 0 | 0 | Negated
denies numbness | 0 | 0 | Negated
denies tingling | 0 | 0 | Negated
denies weakness of the lower extremities | 0 | 0 | Negated
prominent holosystolic murmur at the apex | 0 | 0 | Factual
petechial rash scattered on the abdomen | 0 | 0 | Factual
petechial rash scattered on the palms | 0 | 0 | Factual
petechial rash scattered on the soles of the feet | 0 | 0 | Factual
encephalopathy | 0 | 0 | Factual
facial droop | 0 | 0 | Factual
slurred speech | 0 | 0 | Factual
admitted to the intensive care unit | 0 | 0 | Factual
started on empiric antibiotic treatment with vancomycin | 0 | 72 | Factual
started on empiric antibiotic treatment with meropenem | 0 | 72 | Factual
became unresponsive to voice | 24 | 24 | Factual
minimally responsive to pain | 24 | 24 | Factual
left hemi-neglect | 24 | 24 | Factual
right gaze deviation | 24 | 24 | Factual
Glasgow Coma Scale (GCS) was 6 | 24 | 24 | Factual
intubated for airway protection | 24 | 24 | Factual
leukocytosis of 24.7 × 10^9/L | 0 | 0 | Factual
87.6% neutrophils | 0 | 0 | Factual
platelet count of 17 × 10^9/L | 0 | 0 | Factual
declined a HIV test | 0 | 0 | Factual
innumerable acute to subacute embolic infarcts in both cerebral and cerebellar hemispheres | 0 | 0 | Factual
proximal right internal carotid artery T-shaped acute thrombus | 0 | 0 | Factual
occlusion of the right middle cerebral artery | 0 | 0 | Factual
subarachnoid hemorrhage in the right parietal region | 0 | 0 | Factual
subarachnoid hemorrhage around the posterior aspect of the midbrain | 0 | 0 | Factual
echo densities on the tricuspid valve | 0 | 0 | Factual
echo densities on the aortic valve | 0 | 0 | Factual
echo densities on the mitral valve | 0 | 0 | Factual
blood culture grew S. marcescens | 0 | 0 | Factual
antibiotic changed to cefepime | 72 | 72 | Factual
cardiothoracic surgery consulted | 72 | 72 | Factual
poor candidate for surgery | 72 | 72 | Factual
neurological status continued to deteriorate | 72 | 144 | Factual
no cough or gag reflex | 144 | 144 | Factual
pupils were fixed and mid-dilated | 144 | 144 | Factual
withdrew care | 144 | 144 | Factual
discharged to hospice care | 144 | 144 | Factual