43 years old | 0
male | 0
admitted to the hospital | 0
uncontrolled diabetes mellitus | -336
chronic kidney disease | -336
infected surgical wound | -336
intangible trauma | -336
Ray's amputation | -336
pus in wound | -336
cellulitis | -336
purulent discharge | -336
decreased urination | 0
Foley catheter insertion | 0
leukocytes 17.1 thousands/μL | 0
neutrophils 15.5 thousands/μL | 0
lymphocytes 1.1 thousands/μL | 0
hemoglobin 7.9 g/dL | 0
hematocrit 26.9% | 0
platelets 100 units/μL | 0
fasting blood sugar 175 mg/dL | 0
creatinine 3.5 mg/dL | 0
blood urea nitrogen 189 mg/dL | 0
bilirubin, total 3.7 mg/dL | 0
pH 7.34 | 0
PCO2 30.2 mmHg | 0
HCO3 16.6 Mmol/L | 0
admitted to ICU | 0
vancomycin 1 g/bid | 0
piperacillin/tazobactam 3.376 g/QID | 0
imipenem 500 mg/BID | 0
wound irrigation | 0
sepsis | 0
fever (38.5°C) | 168
systolic hypotension | 168
confusion | 168
leukocytes 12.7 ×10³ | 168
hemoglobin 6.9 g/dL | 168
thrombocytes 39,000/μL | 168
creatinine increased | 168
Guillotine ankle amputation | 168
sepsis control | 240
no purulent discharge | 240
necrotic ulcer | 240
IV injection site involvement | 240
extensive debridement | 240
pathology evaluation | 240
CM diagnosis | 240
amphotericin B 300 mg daily | 240
pulseless radial and ulnar arteries | 288
occlusive clot formation | 288
acute deep vein thrombosis | 288
surgical embolectomy | 288
sepsis persistence | 288
multi-organ failure | 288
death | 288
