46 years old | 0
    African American | 0
    man | 0
    uncontrolled diabetes mellitus | 0
    hypertension | 0
    chronic kidney disease | 0
    polysubstance abuse | 0
    alcohol abuse | 0
    tobacco abuse | 0
    marijuana abuse | 0
    cocaine abuse | 0
    confusion | 0
    difficulty speaking | 0
    temperature 37.6°C (99.7°F) | 0
    blood pressure 154/93 mm Hg | 0
    oriented to self | 0
    expressive (Broca’s) aphasia | 0
    non-fluent speech | 0
    impaired naming | 0
    impaired repetition | 0
    able to follow two-step commands | 0
    good comprehension | 0
    dysarthria | 0
    right-sided hemiparesis | 0
    leukocytosis 12.86 × 10³/μL | 0
    computer tomography left thalamic mass 3.1 cm | 0
    5 mm rightward midline shift | 0
    magnetic resonance imaging confirmed | 0
    admitted to neurological intensive care unit | 0
    empiric intravenous vancomycin | 0
    empiric intravenous meropenem | 0
    stereotactic aspiration | 0
    purulent material | 0
    Gram positive cocci in chains | 0
    Streptococcus anginosus culture | 0
    negative blood cultures | 0
    transthoracic echocardiogram negative for valvular vegetations | 0
    computer tomography sigmoid colitis | 0
    deferred endoscopic evaluation | 0
    antibiotic switched to ceftriaxone | 0
    left against medical advice | 360
    neurosurgery outpatient wound assessment | 720
    persistence of hemiparesis | 720
    no documentation regarding aphasia | 720
    subcortical aphasia | 0
    thalamic brain abscess | 0
    area of sigmoid colitis | 0
    encephalopathy | 0
    contralateral hemiparesis | 0
    expressive aphasia | 0
    deep-seated abscess | 0
    vasogenic edema | 0
    intravenous antimicrobials | 0
    resolution of abscesses | 0
    intraventricular rupture risk | 0
    permanent neurological damage risk | 0
    mortality risk | 0
    morbidity risk | 0
    follow up imaging | 720
    therapeutic end point | 720
    resolution of disease | 720

    46 years old | 0  
African American | 0  
man | 0  
uncontrolled diabetes mellitus | 0  
hypertension |5 0  
chronic kidney disease | 0  
polysubstance abuse | 0  
alcohol abuse | 0  
tobacco abuse | 0  
marijuana abuse | 0  
cocaine abuse | 0  
confusion | 0  
difficulty speaking | 0  
temperature 37.6°C (99.7°F) | 0  
blood pressure 154/93 mm Hg | 0  
oriented to self | 0  
expressive (Broca’s) aphasia | 0  
non-fluent speech | 0  
impaired naming | 0  
impaired repetition | 0  
able to follow two-step commands | 0  
good comprehension | 0  
dysarthria | 0  
right-sided hemiparesis | 0  
leukocytosis 12.86 × 10³/μL | 0  
computer tomography left thalamic mass 3.1 cm | 0  
5 mm rightward midline shift | 0  
magnetic resonance imaging confirmed | 0  
admitted to neurological intensive care unit | 0  
empiric intravenous vancomycin | 0  
empiric intravenous meropenem | 0  
stereotactic aspiration | 0  
purulent material | 0  
Gram positive cocci in chains | 0  
Streptococcus anginosus culture | 0  
negative blood cultures | 0  
transthoracic echocardiogram negative for valvular vegetations | 0  
computer tomography sigmoid colitis | 0  
deferred endoscopic evaluation | 0  
antibiotic switched to ceftriaxone | 0  
left against medical advice | 360  
neurosurgery outpatient wound assessment | 720  
persistence of hemiparesis | 720  
no documentation regarding aphasia | 720  
subcortical aphasia | 0  
thalamic brain abscess | 0  
area of sigmoid colitis | 0  
encephalopathy | 0  
contralateral hemiparesis | 0  
expressive aphasia | 0  
deep-seated abscess | 0  
vasogenic edema | 0  
intravenous antimicrobials | 0  
resolution of abscesses | 0  
intraventricular rupture risk | 0  
permanent neurological damage risk | 0  
mortality risk | 0  
morbidity risk | 0  
follow up imaging | 720  
therapeutic end point | 720  
resolution of disease | 720