62 years old | 0
male | 0
admitted to the hospital | 0
dyspnea | -72
intermittent chest pain | -72
end-stage renal disease | -672
peritoneal dialysis | -672
type 2 diabetes mellitus | -672
aortic stenosis | -672
transcatheter aortic valve implantation (TAVI) | -336
COVID-19 | -24
anemic | -24
progressively hypoxic | -24
intubated | -24
transferred to a tertiary care facility | -24
treated for presumed cytokine storm | -24
hypotension | 0
cardiology consultation | 0
evaluation of aortic valve prosthesis | 0
POCUS performed | 0
large pericardial effusion | 0
cardiac tamponade | 0
advanced cardiac life support initiated | 0
pericardiocentesis performed | 0
60 mL of serous fluid aspirated | 0
return of spontaneous circulation | 0
repeat POCUS performed | 0
decrease in effusion size | 0
expansion of the heart | 0
guide wire advanced | 0
pigtail placed | 0
650 mL of fluid drained | 0
repeat echo performed | 0
resolution of pericardial effusion | 0
normal LV function | 0
discharged | 24