female | 0
infant | 0
born | 0
38 weeks of gestation | 0
cesarean section | 0
first-degree consanguineous marriage | -672
mother 29 years old | -672
no history of radiation exposure | -672
no drug intake during pregnancy | -672
no similar conditions in family | -672
referred to neonatal intensive care unit | 20
suspected duodenal atresia | 20
weight 2400g | 20
length 55cm | 20
head circumference 35cm | 20
stable vital signs | 20
afebrile | 20
heart rate 130/minute | 20
respiratory rate 55/minute | 20
oxygen saturation 95-96% | 20
normal blood investigations | 20
normal platelets | 20
deformity of left upper limb | 20
radial flexion | 20
partial syndactyly | 20
complete radial aplasia | 20
abnormal flexion of wrist | 20
no other osseous anomalies | 20
soft abdomen | 20
passing stool | 20
nil per os | 20
dilated stomach | 20
residual gastric greenish aspirate | 20
suspected duodenal web | 20
laparotomy | 48
annular pancreas | 48
obstructing duodenum | 48
dilated stomach and duodenum | 48
normal liver | 48
patent hepatic veins | 48
gall bladder | 48
normal kidneys | 48
no ascites | 48
no spleen | 48
Howell-Jolly bodies | 48
absence of spleen | 48
asplenia syndrome | 48
standard spleen and liver scan | 48
normal liver location | 48
no spleen visualized | 48
levocardia | 48
complex congenital heart disease | 48
single atrium | 48
single ventricle | 48
single AV valve | 48
dextro-transposition of great arteries | 48
moderate pulmonary valve stenosis | 48
small patent ductus arteriosus | 48
normal head ultrasound | 48
small focus of increased parenchymal echogenicity | 48
persistent late-onset staphylococcus sepsis | 504
prolonged antibiotic treatment | 504
full feeding | 504
extubated to nCPAP | 504
oxygen requirement 30% | 504
prophylactic antibiotic therapy | 504
anti-heart failure medications | 504
follow-up with cardiology | 504
follow-up with orthopedic | 504
follow-up with plastic surgeons | 504
accepted for further management | 504
discharged | 720