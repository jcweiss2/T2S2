58 years old | 0
male | 0
admitted to the hospital | 0
6-month headache | -4320
progressive right hemiparesis | -4320
hyperreflexia | 0
positive right Babinski reflex | 0
computed tomography scan | 0
left thalamic lesion | 0
ring-enhancement pattern | 0
leukocytosis | 0
negative detection of anti-HIV antibodies | 0
VITEK MS analysis | 0
N. beijingensis infection | 0
triple antibiotic therapy | 0
meropenem | 0
trimethoprim/sulfamethoxazole | 0
amikacin | 0
ventriculostomy system | 0
Ommaya reservoir | 0
blood and cerebrospinal fluid cultures | 0
thoracoabdominal CT scan | 0
no mass or solid organ lesion | 0
transthoracic and transesophageal echocardiograms | 0
no endocarditis | 0
clinical improvement | 168
seizure episode | 168
anisocoria | 168
emergency CT scan | 168
orotracheal intubation | 168
severe swelling | 168
increase in abscess size | 168
supratentorial ventriculomegaly | 168
cisternal obstruction | 168
emergency Ommaya puncture | 168
turbid-yellow liquid | 168
abscess drained | 168
capsule partially resected | 168
contralateral ventriculostomy system | 168
systemic inflammatory response syndrome | 192
Pseudomonas aeruginosa | 192
Klebsiella pneumoniae | 192
tracheitis | 192
vancomycin | 192
fever | 192
tachycardia | 192
multilobed opacities | 192
gram-positive bacilli | 192
septic shock | 192
pulmonary foci | 192
multiple antibiotic regimen | 192
vasoactive support | 216
anticonvulsive management | 216
myoclonic movements | 216
death | 336
intraoperative sample | -4320
N. beijingensis | -4320
hsp65 | 0
16S-23S rRNA gene intergenic spacer | 0
genotyping | 0
PCR products | 0
Sanger method | 0
MEGA-X | 0
NCBI nucleotide collection | 0