37 years old | 0
female | 0
occipital craniectomy | 0
general anesthesia | 0
severe macroglossia | 0
extubation | 0
tracheostomy | 0
posterior occipital lesion | 0
low-grade glioma | 0
pilocytic features | 0
occipital craniotomy | 0
supratentorial approach | 0
tumor debulking | 0
ASA II | 0
unremarkable physical exam | 0
no allergies | 0
left parietal craniotomy | -144000
partial tumor excision | -144000
chemotherapy | -144000
radiotherapy | -144000
increased intracranial pressure | -144000
EVD insertion | -144000
recurrence of brain tumor | -105120
right occipital craniotomy | -105120
metastatic sub-thalamic brain tumor | -96000
blurred vision | -96000
navigation-assisted tumor debulking | -96000
surgical procedure (10 hours) | 0
sitting position | 0
minimal head flexion | 0
throat pack insertion | 0
invasive monitoring | 0
left radial arterial line | 0
right subclavian central line | 0
propofol induction | 0
fentanyl induction | 0
cisatracurium muscle relaxation | 0
cuffed ETT (7.5 mm) | 0
Cormack-Lehane grade 1 view | 0
mechanical ventilation | 0
isoflurane maintenance | 0
cisatracurium infusion (8 mg/hour) | 0
remifentanil infusion |5| 0
Ringer lactate (3.5 liters) | 0
PRBCs transfusion | 0
adequate urine output | 0
stable vital signs | 0
systolic blood pressure (~100 mmHg) | 0
PaCO2 (~33 mmHg) | 0
oxygen saturation (99%) | 0
residual muscle paralysis reversal | 0
neostigmine | 0
atropine | 0
throat pack removal | 0
spontaneous breathing | 0
tidal volume (800–850 mL) | 0
respiratory rate (10–12 breaths/min) | 0
neurological exam (left-sided weakness) | 0
neurosurgery team informed | 0
slipped head dressing | 0
gradual decrease in tidal volume | 0
rapid tongue size increase | 0
O2 saturation decreased (early 90s%) | 0
manual mask ventilation | 0
high resistance | 0
foreign body suspicion | 0
oropharynx checked by laryngoscope | 0
enlarged tongue | 0
edematous soft palate | 0
Cormack-Lehane grade 4 | 0
difficult intubation | 0
mask ventilation harder | 0
inspiratory stridor | 0
O2 saturation dropped (80s%) | 0
call for help | 0
O2 saturation maintained (93–94%) | 0
no fiber-optic trial | 0
surgery team consulted for tracheostomy | 0
bag-mask ventilation difficulty | 0
tracheostomy without complications | 0
ICU transfer | 0
propofol sedation | 0
remifentanil sedation | 0
cefuroxime | 0
vancomycin | 0
levofloxacin | 0
dexamethasone | 0
antihistamine | 0
enteral feeding | 0
nasogastric tube | 0
chest physiotherapy | 0
macroglossia (Figure 1A) | 0
increased tongue and neck swelling (2 days later) | 48
mouth gag application | 48
MRA ordered | 48
MRA not done | 48
increased WBC count (5 days later) | 120
septic work-up | 120
gram-negative bacilli | 120
tongue size increase (9 days later) | 216
ulcerations on tongue surface | 216
sepsis (16 days later) | 384
multi-organ failure | 384
asystole | 384
death | 384
