37 years old | 0
    primigravida | 0
    twin gestation | 0
    admitted | 0
    epigastric discomfort | 0
    abdominal pain | 0
    malaise | 0
    vomiting | 0
    hypertension | 0
    third trimester | 0
    alpha methyldopa | 0
    heart rate 102/min | 0
    blood pressure 170/90 mm Hg | 0
    icterus | 24
    fetal heart sounds | 0
    ultra sonography fatty liver | 0
    ultra sonography twin pregnancy | 0
    haemoglobin 10.7 g% | 0
    total count 10,700/mm3 | 0
    platelets 2.6 lakhs | 0
    urea 11 mg/dl | 0
    creatinine 1.4 mg/dl | 0
    uric acid 5.3 mg/dl | 0
    lactate dehydrogenase 442 U/L | 0
    peripheral smear negative for haemolysis | 0
    Hepatitis B surface antigen negative | 0
    Hepatitis C virus negative | 0
    Human immunodeficiency virus negative | 0
    prothrombin time test 48 s control 14 s | 0
    International Normalised Ratio 4.0 | 0
    total bilirubin 7.8 mg/dl | 0
    direct bilirubin 4.0 mg/dl | 0
    serum glutamic oxaloacetic transaminase 316 U/L | 0
    serum glutamic-pyruvic transaminase 313 U/L | 0
    alkaline phosphatase 974 | 0
    total protein 5.3 U/L | 0
    albumin 2.8 U/L | 0
    globulin 2.5 U/L | 0
    plasma ammonia 93 meq/d | 0
    urine albumin++ | 0
    cardiotocography fetal distress | 0
    pre-eclampsia | 0
    acute fatty liver of pregnancy | 0
    emergency caesarean section | 0
    vitamin K | 0
    fresh frozen plasma | 0
    general anesthesia | 0
    induction by rapid sequence | 0
    thiopentone | 0
    suxamethonium | 0
    trachea intubated | 0
    endotracheal tube size seven | 0
    oxygen | 0
    nitrous oxide | 0
    sevoflurane | 0
    fentanyl | 0
    atracurium | 0
    mannitol | 0
    albumin transfused | 0
    twin babies delivered | 0
    extubation | 0
    recovery uneventful | 0
    cryoprecipitate | 0
    fresh frozen plasma transfused | 0
    broad spectrum antibiotics started | 0
    magnesium sulphate continued at 2 g/h | 0
    serum magnesium levels monitored | 0
    liver function deteriorated further | 72
    tonic clonic convulsions | 96
    respiratory distress | 96
    chest X-ray acute respiratory distress syndrome | 96
    mechanical ventilation initiated | 96
    antibiotic changed to tobramycin | 96
    computed tomography scan brain normal | 96
    electroencephalography normal | 96
    repeat ultra sound scan ascites | 96
    hyperechoic features haemorrhagic ascites | 96
    coagulopathy | 96
    no gall stones | 96
    no dilatation of biliary tract | 96
    central venous pressure maintained 8-12 mm Hg | 96
    weaned off | 168
    non-invasive ventilation continued | 168
    hepatic function gradually improved | 168
    viral markers negative | 168
    coagulopathy corrected | 480
    patient gradually improved | 480
    shifted out from post-operative intensive care unit | 480