72 years old | 0
male | 0
dermatomyositis | -480
pancytopenic | -120
methotrexate therapy | -120
aplastic anemia | -120
bone marrow biopsies | -120
hypocellularity | -120
neutropenic fever | -24
hospitalization | -24
ATG therapy | 0
ID skin test | 0
wheal and flare reaction | 0
prednisone | 0
total white blood cell count | 0
lymphocytes | 0
epicutaneous skin test | 120
histamine control | 120
saline control | 120
desensitization | 120
informed consent | 120
desensitization regimen | 120
intensive care unit | 120
diphenhydramine | 120
ranitidine | 120
acetaminophen | 120
methylprednisolone | 120
ATG desensitization | 120
increasing dilutions of ATG | 120
premedication | 120
rescue medications | 120
full therapeutic dosing | 144
fungal septicemia | 672
death | 672
ID skin test positive | 0
epicutaneous skin test negative | 120
anaphylaxis | -120
desensitization protocol | 120
ATG hypersensitivity | 0
type I hypersensitivity | 0
epicutaneous skin testing | 120
ID skin testing | 0
specific IgE | 120
false positive ID skin test | 120
localized side effects | 120
systemic side effects | 120
successful desensitizations | 120
ATG package insert | 0
epicutaneous testing | 120
ID testing | 0
drug desensitization | 120
anaphylaxis management | 120