74 years old | 0
male | 0
admitted to the hospital | 0
head trauma | -24
fall | -24
bruises on arms and legs | -24
dementia | 0
Glasgow Coma Scale 13/15 | 0
heart rate 94 beats per minute | 0
blood pressure 149/75 mmHg | 0
temperature 37.9°C | 0
abrasion wound on head | 0
bruises on chest and upper abdomen | 0
severe tenderness in right lower leg | 0
MMT four-fifths in right lower leg | 0
hemoglobin 13.5 mg/dL | 0
leukocyte count 19,200 cells/μL | 0
neutrophil count 15,398 cells/μL | 0
urea 25 mmol/L | 0
creatinine 0.76 mg/dL | 0
potassium 3.8 mmol/L | 0
sodium 141 mmol/L | 0
chloride 108 mmol/L | 0
creatine kinase 20,518 IU/L | 0
C-reactive protein 13.43 mg/dL | 0
tetanus vaccine administered | 0
intravenous tazobactam/piperacillin hydrate | 0
no fractures on upper limbs, lower limbs, or pelvis | 0
SAH | 0
acute subdural hematoma | 0
hypodense lesions in bilateral parietooccipital areas | 0
no fractures of cranial bones | 0
no abnormalities in lung and abdominal CT | 0
no carotid stenosis | 0
no brain aneurysm | 0
no vasospasm | 0
cortical and subcortical altered intensities in bilateral parietooccipital areas | 0
hyperintense regions on T2WI | 0
hyperintense regions on FLAIR | 0
hyperintense regions on DWI | 0
hyperintense regions on ADC | 0
normal spinal cord MR imaging | 0
ascending weakness in extremities | 48
bulbar weakness | 48
complete quadriplegia | 288
bulbar palsy | 288
weakness of respiratory muscles | 288
lower oxygen saturation | 288
respiratory intubation | 288
mechanical ventilation | 288
absent DTR | 288
unclear sensory loss | 288
possible GBS | 288
IVIg administered | 288
leukocyte count 12,700 cells/μL | 288
C-reactive protein 3.50 mg/dL | 288
creatine kinase within normal limits | 288
no anti-GM1 antibodies | 288
no anti-GQ1b antibodies | 288
negative blood cultures | 288
negative CSF cultures | 288
no Epstein–Barr virus detected | 288
no herpes simplex detected | 288
no cytomegalovirus detected | 288
CSF protein 92 mg/dL | 288
CSF cell count 8/mmc | 288
no electrophysiological analysis | 288
increased signals on T2WI | 288
increased signals on FLAIR | 288
increased signals on DWI | 288
increased signals on ADC | 288
extubated | 576
improved MMTs of limbs | 576
brisk DTR | 576
disappearance of T2WI hyperintensities | 576
disappearance of FLAIR hyperintensities | 576
disappearance of DWI hyperintensities | 576
disappearance of ADC hyperintensities | 576
sent to rehabilitation hospital | 1320
antibiotic-resistant pyrexia | 72
neurogenic fever | 72
no respiratory symptoms | 0
no abdominal symptoms | 0
no infection findings | 0
no electrolyte disturbance | 0
no botulism | 0
no myasthenia gravis | 0
no periodic paralysis | 0
no poliomyelitis | 0
rhabdomyolysis | 0
PRES diagnosis | 576
possible GBS diagnosis | 288
resolution of PRES | 576
resolution of GBS | 576
