67 years old | 0
male | 0
admitted to the hospital | 0
fever | 0
lethargy | 0
tachycardia | 0
tachypnea | 0
hypotension | 0
aorto-bi-iliac graft replacement | -8760
Abdominal Aortic Aneurysm (AAA) | -8760
paraplegia | -8760
graft leaking | -8760
embolization | -8760
intubation | 0
transferred to the medical critical care unit | 0
White blood cell count 17,000/μL | 0
Hemoglobin 9.6 g/dL | 0
platelet count 300,000/μL | 0
BUN 66 mg/dL | 0
Cr 2.1 mg/dL | 0
minimal elevation of troponin | 0
normal level of electrolytes | 0
severe sepsis | 0
septic shock | 0
vancomycin | 0
Meropenem | 0
Eggerthella lenta | 0
Escherichia coli Extended-spectrum beta-lactamase (ESBL) | 0
Enterococcus Faecalis | 0
transesophageal echocardiogram | 0
no vegetation | 0
Abdominal computed tomography (C.T.) | 0
inflammatory changes around aorto-bi-iliac graft | 0
no aortoenteric fistula | 0
Indium-111 WBC scan | 24
abnormally increased activity in the mid to lower abdomen | 24
vascular surgery evaluation | 0
conservative strategy | 0
IV antibiotics | 0
vancomycin (1 g daily) | 0
Meropenem (1 g twice a day) | 0
spiking of fever | 168
unable to be weaned from mechanical ventilation | 168
repeat blood culture | 168
Tigecycline (50 mg twice a day) | 168
repeat blood cultures were negative | 170
discharged home | 336
long term antibiotic therapy | 336
close control of inflammation markers | 336