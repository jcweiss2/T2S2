49 years old | 0
male | 0
African American | 0
morbidly obese | 0
end-stage renal disease | 0
peritoneal dialysis | 0
hypertension | 0
nausea | -96
nonbilious nonbloody emesis | -96
severe diffuse abdominal pain | -96
reported symptoms to outpatient PD nurse | -48
cloudy white fluid | -48
peritoneal fluid and culture sent for evaluation | -48
started on intraperitoneal cefazolin | -48
started on intraperitoneal ceftazidime | -48
fever | -24
temperature 101.5 °F | -24
admitted to hospital | 0
afebrile | 0
blood pressure 95/72 mmHg | 0
heart rate 88 bpm | 0
respiratory rate 20 breaths/min | 0
acute distress secondary to abdominal pain | 0
distended abdomen | 0
tender to light palpation | 0
positive fluid wave | 0
dull to percussion | 0
leukocytosis | 0
potassium 3.3 mmol/L | 0
anion gap 25 | 0
peritoneal fluid total white blood cell count 93 557 | -48
neutrophil predominance 80% | -48
Acinetobacter pittii identified | 24
started on intraperitoneal ceftazidime and gentamicin | 24
susceptibilities returned | 48
sensitive to ceftazidime | 48
blood culture results showed no growth | 120
continued on intraperitoneal ceftazidime | 120
treatment extended to 28 days | 336
readmitted to hospital | 816
fever | 816
abdominal pain | 816
peritoneal fluid cell count elevated | 816
cultures growing Acinetobacter pittii | 816
started on vancomycin and gentamicin | 816
started on intravenous ceftazidime | 816
PD catheter removed | 840
hemodialysis initiated | 840
discharged with ciprofloxacin | 864
asymptomatic upon completion of therapy | 888