69 years old | 0
male | 0
admitted to the ICU | -336
pneumonia | -336
mitral valve surgery | -336
severe sepsis | -336
treated with high doses of vasopressors | -336
required continuous hemodialysis | -336
invasive ventilator support | -336
remifentanil infusion | -336
decannulated | -168
hyperactive delirium | -168
confusion | -168
paranoia | -168
hallucinations | -168
agitation | -168
non-pharmacological treatment | -168
early mobility | -168
sleep-wake cycle preservation | -168
olanzapine prescribed | -168
10 mg olanzapine orally | -168
dosage changed to twice daily | -24
fourth dose of olanzapine | 0
hypotensive | 0.5
blood pressure 70/40 mmHg | 0.5
heart rate 90 beats per min | 0.5
nonresponsive | 2
Glasgow coma scale score 7 | 2
pinpoint pupils | 2
airway maintained | 2
respiratory rate elevated | 2
arterial blood gas showed normal pO2 | 2
low pCO2 | 2
blood sugar level slightly elevated | 2
norepinephrine infusion started | 2
Glasgow coma scale score remained at 7 | 2
naloxone administered | 2.25
no effect | 2.25
flumazenil administered | 2.5
symptoms reversed | 2.5
pupils dilated back to normal | 2.5
zolpidem administered | -12
ipratropium inhalations | -12
dalteparin administered | 0
esomeprazole administered | 0
macrogol administered | 0
meropenem administered | 0
micafungin administered | 0
mirtazapine administered | 0
nicotine transdermal patch | 0
paracetamol administered | 0
potassium citrate administered | 0
pregabalin administered | 0
salbutamol inhalation | 0
zopiclone administered | -2