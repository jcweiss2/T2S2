43 years old | 0
    male | 0
    diabetes mellitus | 0
    hypertension | 0
    recovered from COVID-19 | -72
    blurred vision on left eye field | -72
    impaired vision on left eye field | -72
    retro-orbital pain | -72
    headache | -72
    transient relief of symptoms | -72
    symptoms recurred | -72
    visual acuity 6/36 left eye | 0
    visual acuity 6/6 right eye | 0
    impaired abduction left eye | 0
    impaired upward movement left eye | 0
    impaired vision left eye | 0
    relative afferent pupillary defect left eye | 0
    brisk reflex right eye | 0
    blurred disc margin left eye | 0
    flat retina both eyes | 0
    hematocrit 42% | 0
    white blood cell count 14500/uL | 0
    neutrophils 95% | 0
    lymphocytes 5% | 0
    erythrocytes sedimentation rate 31 mm/h | 0
    optic neuritis | -72
    heterogeneously enhancing lesion left orbital apex | 0
    lesion encasing left optic nerve | 0
    lesion compressing left optic nerve | 0
    focal asymmetric enhancement left cavernous sinus | 0
    heterogeneously enhancing soft tissue left orbital apex | 0
    widening of canal | 0
    mild extension into sphenoid sinus | 0
    excision biopsy left orbital apex lesion | 0
    yellowish-white tissue | 0
    purulent discharge | 0
    aspergillosis | 0
    orbital apex syndrome | 0
    IV methylprednisolone for 3 days | -72
    oral prednisolone 60 mg for 2 days | -72
    tapered prednisolone for 1 month | -72
    repeat MRI performed | -72
    no evidence of lesion | -72
    treated again for optic neuritis | -72
    symptoms relief transiently | -72
    pain recurred | -72
    vision impairment recurred | -72
    no longer perceived light OD | -72
    another course of prednisolone | -72
    orbital MRI performed | -72
    paranasal CT scan performed | -72
    denied diplopia | 0
    denied scalp tenderness | 0
    denied weight loss | 0
    denied jaw claudication | 0
    
    <|eot_id|>
