83 years old | 0
male | 0
prostatic cancer | -105120
diabetes mellitus | 0
hypertension | 0
hyperuricemia | 0
lower back pain (gradually progressive) | -1176
admitted to the emergency room | 0
compression fracture of L2 vertebra | -840
painkillers | -840
diagnosed with prostatic cancer | -105120
hormones | -105120
radiation | -105120
treated for diabetes mellitus | 0
treated for hypertension | 0
treated for hyperuricemia |%0
heart rate 140 beats/min | 0
respiratory rate 39 breaths/min | 0
percutaneous arterial oxygen saturation 89% | 0
oxygen therapy via nasal cannula at 2 L/min | 0
lower back pain | 0
tenderness in left thigh | 0
stabbing pain in left thigh | 0
erythematous rash in left thigh | 0
white blood cell count 30,600 cells/mm3 | 0
neutrophils 92.9% | 0
hemoglobin 10.9 g/dL | 0
creatinine 2.48 mg/dL | 0
C-reactive protein 42.72 mg/dL | 0
procalcitonin 29.69 ng/mL | 0
glucose level 156 mg/dL | 0
glycated hemoglobin 6.1% | 0
computed tomography scan | 0
massive pleural effusion in left thoracic cavity | 0
fluid retention in left iliopsoas muscle | 0
air extending to lower limb | 0
inflammation in retroperitoneal cavity | 0
diffuse low-density region in front of lumbar vertebrae | 0
lumbar vertebral infection | 0
Sequential Organ Failure Assessment (SOFA) score 6 | 0
rapid infusion | 0
pressor agents | 0
intravenous meropenem 1 g | 0
thoracotomy tube insertion | 0
drain pleural effusion | 0
exudative effusion | 0
neutrophil count 25,000 cells/μL | 0
abscess in left thigh incised | 0
abscess drained | 0
catheter inserted into retroperitoneal cavity | 0
chocolate-colored pus | 0
foul-smelling pus | 0
admitted to intensive care unit | 0
continuous hemodiafiltration | 0
ventilator control | 0
sepsis management | 0
meropenem 2 g daily | 0
clindamycin 1200 mg daily | 0
died of multiple organ failure | 72
necrotizing fasciitis | 72
myositis | 72
neutrophil infiltration | 72
gram-positive bacteria | 72
anaerobic culture of pleural effusion positive | 96
blood culture needed more few days | 96
Parvimonas micra identified | 96
16S ribosomal RNA match 99.9% | 96
P. micra identified in blood | 96
P. micra identified in pleural fluid | 96
P. micra identified in pus | 96
