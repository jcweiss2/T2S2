62 years old | 0
male | 0
admitted to the hospital | 0
febrile neutropenia | 0
dry cough | 0
dyspnea | 0
autologous bone marrow transplant | -384
mantle cell lymphoma | -384
chest CT | 0
diffuse tracheobronchial thickening | 0
densification of the adjacent mediastinal fat | 0
empirical antibiotic therapy | 0
amphotericin B | 0
follow-up CT | 24
persistence of cough | 24
hemoptysis | 24
worsening of the imaging findings | 736
greater tracheal and bronchial walls thickening | 736
increased densification of the adjacent mediastinal fat | 736
laryngotracheobronchoscopy | 1008
whitish plaques | 1008
friable mucosa | 1008
segmental ostial obstruction | 1008
bronchoalveolar lavage | 1008
endobronchial biopsy | 1008
bifurcated hyphae | 1010
Grocott method | 1010
Aspergillus sp | 1010
disease progression | 1010
bronchoalveolar lavage culture | 1010
positive for Aspergillus sp | 1010
discharged | 1012
oral voriconazol | 1014
abdominal pain | 1016
diarrhea | 1016
hypotension | 1016
febrile peak | 1016
septic shock | 1016
intensive care unit | 1016
death | 1019