40 years old | 0
female | 0
liver transplantation | -304
cirrhosis | -304
nonalcoholic steatohepatitis | -304
hypertrophic cardiomyopathy | -1096
myomectomy | -1096
hypothyroidism | -304
Type II diabetes mellitus | -304
chronic kidney disease | -304
tacrolimus | -304
mycophenolic acid | -304
prednisone | -304
possible tacrolimus-related posterior reversible encephalopathy syndrome | -156
everolimus-based therapy | -156
liver biopsy | -120
severe acute cellular rejection | -120
high-dose steroids | -120
thymoglobulin | -120
cyclosporine | -120
admitted to Intensive Care Unit | 0
adult respiratory distress syndrome | 0
septic shock | 0
Legionella pneumophila pneumonia | 0
respiratory failure | 0
failed extubation | 0
ventilatory support | 0
acute on chronic renal failure | 0
CRRT | 0
propofol | 0
heparin infusion | 0
activated partial thromboplastin time | 0
right radial artery thrombus | 0
CRRT filter clotting | 312
elevated triglycerides | 312
discontinuation of propofol | 312
filter and circuits changed | 312
adjunctive therapy with intravenous insulin | 312
heparin | 312
therapeutic plasma exchange | 318
rising serum potassium | 318
serum bicarbonate | 318
pH | 318
emergent therapeutic plasma exchange | 318
CRRT resumed | 324
new filter | 324
acid-base balance normalized | 324
electrolytes normalized | 324
elevated TG levels | 384
increasing serum lipase levels | 384
abdominal pain | 384
concern for pancreatitis | 384
additional TPE sessions | 384
TG decreased | 384
oral fibrate | 384
fish oil | 384
combined liver-kidney transplant | 1344
propofol for sedation | 1344
cyclosporine postoperatively | 1344
TGs level normalized | 1344
TGs level remained well-controlled | 1344