64 years old | 0
woman | 0
admitted to the clinic | 0
increasing dyspnoea | -72
edema of lower limbs | -72
elevated NT-proBNP | 0
right axis deviation | 0
right atrial enlargement | 0
carcinoid tumor of terminal ileum | -672
hepatic metastasis | -672
lymphatic metastasis | -672
osseous metastasis | -672
partial ileum resection | -672
somatostatin analogue | -672
tumor staging | -672
laboratory evaluation | -672
partial remission | -672
severe pulmonary stenosis | 0
torrential tricuspid regurgitation | 0
coaptation defect | 0
thickening of valve leaflets | 0
retraction of valve leaflets | 0
surgical valve replacement | 24
uneventful surgery | 24
uneventful initial postoperative course | 24
condition worsened | 48
cardiac complications excluded | 48
carcinoid crises excluded | 48
pneumogenic sepsis | 48
broad-spectrum targeted anti-infective therapy | 48
intensive care measures | 48
therapy-refractory multi-organ failure | 72
death | 72
