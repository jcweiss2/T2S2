34 years old | 0
multipara | 0
admitted to the hospital | 0
low abdominal pain | 0
nausea | 0
vomiting | 0
height 157 cm | 0
weight 67 kg | 0
weight gain during pregnancy 13 kg | 0
parity 1-0-0-1 | 0
no abnormalities in past medical history | 0
blood pressure 120/75 mmHg | 0
heart rate 75 beats/min | 0
respiratory rate 22 times/min | 0
normal chest radiography | 0
ST segment depression | 0
increased troponin-T | 0
normal CK-MB | 0
normal lab test | 0
fetal heart rate 130 beats/min | 0
blood pressure increased to 158/100 mmHg | 1
sinus tachycardia | 1
moderate decline in systolic function | 1
moderate mitral regurgitation | 1
tricuspid regurgitation | 1
pulmonary hypertension | 1
LVEF 39% | 1
LVEDD 5.2 cm | 1
LVESD 4.3 cm | 1
transferred to intensive care | 1
blood pressure 149/100 mmHg | 1
heart rate 110 beats/min | 1
respiration rate 27 times/min | 1
hemoptysis | 4
dyspnea | 4
oxygen provided | 4
severe pulmonary edema | 4
furosemide injected | 4
nitroglycerin injected | 4
oxygen supplied through mask | 4
ABGA | 4
fetal distress anticipated | 4
cesarean section decided | 4
severe dyspnea | 5
orthopnea | 5
hemoptysis | 5
blood pressure 130/98 mmHg | 5
heart rate 128 beats/min | 5
respiratory rate 45 times/min | 5
sinus tachycardia | 5
general anesthesia decided | 5
ECMO installation attempted | 5
ECMO installation failed | 5
ECMO installed under general anesthesia | 5
cesarean section performed | 5
oxygen 10 L/min through mask | 5
nitroglycerin 12 µg/min | 5
monitoring started | 5
catheter inserted | 5
blood pressure 135/98 mmHg | 5
heart rate 130 beats/min | 5
peripheral oxygen saturation 98% | 5
ABGA | 5
induction of anesthesia | 5
thiopental sodium injected | 5
succinylcholine injected | 5
intubation performed | 5
atracurium injected | 5
anesthesia maintained | 5
ventilator set | 5
blood pressure 155/110 mmHg | 5
heart rate 138 beats/min | 5
sinus tachycardia | 5
anesthetic ABGA | 5
ECMO applied | 5
return canula inserted | 5
drainage canula inserted | 5
flow rate maintained | 5
central venous catheter inserted | 5
Swan-Ganz catheter attempted | 5
blood pressure maintained | 5
heart rate maintained | 5
peripheral oxygen saturation maintained | 5
central venous pressure maintained | 5
ABGA | 5
ventilator adjusted | 5
nitroglycerin injected | 5
infant delivered | 10
APGA score 3 and 4 | 10
intubation performed | 10
oxytocin injected | 10
colloid solution administered | 10
blood pressure maintained | 10
heart rate maintained | 10
peripheral oxygen saturation maintained | 10
central venous pressure maintained | 10
ABGA | 10
patient transferred to ICU | 100
ECMO maintained | 100
intubation maintained | 100
blood pressure 90-100 mmHg | 100
heart rate 110 beats/min | 100
peripheral oxygen saturation 100% | 100
ABGA | 100
flow speed of ECMO decreased to 2 L/min | 72
blood pressure 95-120/79-95 mmHg | 72
heart rate 90-110 beats/min | 72
peripheral oxygen saturation 100% | 72
central venous pressure 5-8 mmHg | 72
ABGA | 72
mechanical ventilation maintained | 72
flow speed of ECMO decreased to 1.3 L/min | 96
blood pressure 120-140/90-100 mmHg | 96
heart rate 90-100 beats/min | 96
peripheral oxygen saturation 100% | 96
central venous pressure 4-8 mmHg | 96
ABGA | 96
flow speed of ECMO decreased to 1 L/min | 108
blood pressure maintained | 108
mechanical ventilation maintained | 108
blood pressure 110-140/80-100 mmHg | 120
heart rate 80-100 beats/min | 120
peripheral oxygen saturation 100% | 120
central venous pressure 9 mmHg | 120
ABGA | 120
ECMO removed | 120
blood pressure 94-104/66-70 mmHg | 120
heart rate 100 beats/min | 120
peripheral oxygen saturation 100% | 120
central venous pressure 5-7 mmHg | 120
ABGA | 120
dopamine injected | 120
mechanical ventilation removed | 168
patient transferred to general ward | 168
blood pressure 100-130/65-70 mmHg | 168
heart rate 75-90 beats/min | 168
ABGA | 168
ECG normal | 168
pulmonary edema improved | 168
LVEF 58% | 168
mitral regurgitation slight | 168
infant transferred to neonate ICU | 168
intubation maintained | 168
extubation performed | 192
abdominal sonography normal | 192
brain MRI normal | 192
infant discharged | 264