69 years old | 0
female | 0
hypertension | 0
type 2 diabetes mellitus | 0
hypersensitivity pneumonitis | 0
obesity | 0
gastric band placement | 0
right breast cancer | 0
status post-lumpectomy | 0
admitted to the hospital | 0
chest pain | 0
shortness of breath | 0
diaphoresis | 0
regular heart rate and rhythm | 0
no murmurs or gallops | 0
clear lungs | 0
anterior ST elevation | 0
elevated troponin level | 0
ST-elevation myocardial infarction (STEMI) | 0
aspirin | 0
heparin | 0
statin therapy | 0
cardiac catheterization | 0
percutaneous coronary intervention | 0
100% occlusion of the left anterior descending (LAD) artery | 0
aspiration thrombectomy | 0
dual antiplatelet therapy | 0
left upper quadrant abdominal pain | 24
diaphoretic | 48
short of breath | 48
fever | 48
tachycardic | 48
hypotensive | 48
leukocytosis | 48
splenic infarct | 48
high-grade stenosis of the celiac artery | 48
mild thickening of the splenic flexure | 48
transthoracic echocardiography | 48
ejection fraction of 40% | 48
apical and mid/anteroseptal wall hypokinesia | 48
trace pericardial effusion | 48
no significant valvular pathology | 48
cardiogenic shock | 48
milrinone | 48
Swan-Ganz catheter | 48
blood cultures | 48
cefepime | 48
metronidazole | 48
heparin infusion | 48
CT angiography | 48
no emboli in her lungs | 48
gram-positive cocci in pairs and chains | 72
vancomycin | 72
repeat blood cultures | 72
E. faecalis | 96
ampicillin | 96
gentamicin | 96
penicillin | 96
ceftriaxone | 96
urinalysis | 96
urine culture | 96
trace leukocytes | 120
negative nitrites | 120
no growth | 120
repeat blood cultures | 120
gram-positive cocci in pairs and chains | 120
E. faecalis | 120
worsening bilateral pleural and pericardial effusion | 120
DENOVA scoring system | 144
septic embolization | 144
unknown origin of bacteremia | 144
four positive blood cultures | 144
TEE | 144
large mobile vegetation | 144
mitral valve | 144
mild mitral regurgitation | 144
no mitral stenosis | 144
ejection fraction of 40% | 144
cardiothoracic surgery department | 144
mitral valve replacement | 144
pre-cardiac surgery workup | 168
head CT | 168
small asymptomatic focus of subarachnoid hemorrhage | 168
head MRI | 168
multiple emboli | 168
left frontal lobe | 168
MRI of the left spine | 168
discitis | 168
osteomyelitis | 168
L1/L2 | 168
carotid duplex ultrasonography | 168
<50% stenosis | 168
right internal jugular vein thrombus | 168
heparin infusion withheld | 168
fluid aspirated from the gastric band | 192
clear | 192
no concerning findings | 192
esophagogastroduodenoscopy | 192
gastric mucosal atrophy | 192
no concern for infection | 192
colonoscopy | 192
perforation | 192
rectosigmoid junction | 192
endoscopically closed | 192
suture | 192
hemoclip | 192
hypoxic | 192
tachycardic | 192
abdominal pain | 192
noninvasive positive-pressure ventilation | 192
epinephrine | 192
exploratory laparotomy | 192
no intraperitoneal contamination | 192
air in the mesentery | 192
extraperitoneal perforation of the rectum | 192
end-colostomy | 192
intensive care unit | 192
persistently febrile | 216
peritonitis | 216
cardiothoracic surgery department | 216
mitral valve replacement | 216
stress dose of hydrocortisone | 216
hydrocortisone | 216
vancomycin | 216
piperacillin/tazobactam | 216
no growth | 240
tracheal aspirate | 240
fever | 240
antibiotic regimen | 240
ceftriaxone | 240
ampicillin | 240
ventilator-associated pneumonia | 264
Stenotrophomonas maltophilia | 264
acute kidney injury | 264
inpatient rehabilitation | 264
acute-on-chronic heart failure | 288
cardiogenic versus septic shock | 288
multiorgan failure | 288
died | 288