54 years old | 0
male | 0
obese | 0
admitted to the hospital | 0
positive coronavirus nasopharyngeal swab test | -120
fever | 0
rigors | 0
persistent cough | 0
myalgia | 0
shortness of breath | 0
no chest pain | 0
no palpitation | 0
no hemoptysis | 0
non-smoker | 0
no alcohol use | 0
no history of liver disease | 0
no co-morbidities | 0
temperature of 39.5 °C | 0
low O2 saturation | 0
blood pressure of 140/82 mm Hg | 0
heart rate of 95/min | 0
respiratory rate of 22/min | 0
bibasilar crackles | 0
no pleural rub | 0
no pericardial rub | 0
no deep vein thrombosis | 0
lymphopenia | 0
high CRP | 0
ferritin 1,620 µg/L | 0
elevated LDH | 0
normal clotting | 0
normal liver function | 0
normal renal function | 0
atypical pneumonia screen negative | 0
blood cultures negative | 0
type 1 respiratory failure | 0
bilateral patchy consolidation | 0
COVID-19 pneumonia | 0
O2 therapy | 0
intravenous antibiotics | 0
dexamethasone | 0
remdesivir | 0
high-flow O2 | 0
tocilizumab | 0
discharged | 0
readmitted | 360
extreme fatigue | 360
poor appetite | 360
reduced oral intake | 360
high temperature | 360
heart rate of 132/min | 360
pyrexial at 38.2 °C | 360
hypotensive | 360
blood pressure of 92/52 mm Hg | 360
tachypnea | 360
respiratory rate of 32/min | 360
GCS 14/15 | 360
icterus | 360
peripherally cyanosed | 360
flapping tremors | 360
encephalopathic | 360
distended tender abdomen | 360
severe type 1 respiratory failure | 360
severe metabolic acidosis | 360
acute kidney injury | 360
hyperkalemia | 360
high creatinine | 360
reduced GFR | 360
acute hepatic injury | 360
elevated ALT | 360
elevated AST | 360
bilirubin elevated | 360
amylase elevated | 360
ALP elevated | 360
GGT elevated | 360
hypoalbuminemia | 360
undetectable paracetamol level | 360
coagulopathy | 360
high INR | 360
raised aPTT | 360
high D-dimer | 360
low platelets | 360
CRP elevated | 360
ferritin extremely high | 360
hemodynamic support | 360
respiratory support | 360
central venous catheter | 360
high-flow oxygen | 360
intubation | 360
ventilation | 360
intravenous piperacillin/tazobactam | 360
intravenous fluids | 360
human albumin serum | 360
fresh frozen plasma | 360
dexamethasone | 360
proton pump inhibitors | 360
bicarbonate | 360
CXR | 360
CT of abdomen and pelvis | 360
multiorgan failure | 360
best supportive care | 360
GCS drop | 360
hypotension | 360
cardiac arrest | 360
death | 384
