65 years old | 0
    female | 0
    diabetes mellitus | 0
    systemic arterial hypertension | 0
    transesophageal echocardiography (TEE) | 0
    suspected diagnosis of atrial septal defect | 0
    procedure performed without sedation | 0
    topical anesthesia | 0
    three attempts of procedure | 0
    procedure interrupted | 0
    difficulties in progression of the probe into the esophagus | 0
    retching | 0
    inability to collaborate with exam performance | 0
    neck pain | 0
    oropharyngeal pain | 0
    severe dysphagia | 24
    edema | 48
    hyperemia | 48
    anterior neck surface pain | 48
    weakness | 48
    malaise | 48
    admitted to the hospital | 72
    looked well | 72
    blood pressure 150/100 mmHg | 72
    pulse rate 100 beats per minute | 72
    edema evident on anterior neck surface | 72
    hyperemia evident on anterior neck surface | 72
    subcutaneous emphysema palpable | 72
    oropharynx hyperemia | 72
    computed tomography (CT) scan of the neck | 72
    subcutaneous emphysema in mediastinal space | 72
    subcutaneous emphysema in supraclavicular space | 72
    subcutaneous emphysema in retroesophageal space | 72
    fistula of posterior esophageal wall at C6–C7 level | 72
    upper gastrointestinal endoscopy | 72
    marked vascular congestion | 72
    edema of hypopharynx | 72
    progression to pyriform sinuses | 72
    progression to upper esophageal sphincter | 72
    obstruction hindering examination | 72
    2 cm perforation of esophageal wall | 72
    purulent secretion draining | 72
    remaining endoscopic examination normal | 72
    diagnosis of esophageal injury | 72
    mediastinal involvement | 72
    ceftriaxone initiated | 72
    clindamycin initiated | 72
    cervicotomy carried out | 72
    drainage of pus from upper mediastinum | 72
    drainage of pus from periesophageal space | 72
    septic shock | 72
    norepinephrine required | 72
    mechanical ventilatory support | 72
    intensive care for a week | 168
    clinical status improved | 168
    esophageal fistula remaining | 168