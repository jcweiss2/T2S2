24 years old | 0 | 0 
female | 0 | 0 
pregnancy | -156 | 0 
abdominal pain | -120 | 0 
abdominal distension | -120 | 0 
constipation | -120 | 0 
admitted to the hospital | 0 | 0 
dehydrated | 0 | 0 
hypotension | 0 | 0 
tachycardia | 0 | 0 
tachypnea | 0 | 0 
asymmetrically distended abdomen | 0 | 0 
tenderness all over abdomen | 0 | 0 
empty rectum on digital examination | 0 | 0 
foetal viability assessed | 0 | 0 
vaginal examination | 0 | 0 
elevated white cell count | 0 | 0 
urine analysis clear | 0 | 0 
ultrasound scan of abdomen and pelvis | 0 | 0 
distended bowel loop | 0 | 0 
free fluid in peritoneal cavity | 0 | 0 
single viable foetus | 0 | 0 
abdominal X-ray | 0 | 0 
dilated large bowel | 0 | 0 
abnormal gas pattern | 0 | 0 
coffee bean appearance | 0 | 0 
sigmoid volvulus diagnosed | 0 | 0 
gastroenterology team consulted | 0 | 0 
emergency sigmoidoscopy | 0 | 0 
twisted sigmoid colon | 0 | 0 
obstruction not negotiated | 0 | 0 
foetal distress | 0 | 0 
deceleration in heart rate | 0 | 0 
concomitant caesarean section | 0 | 0 
premature foetus delivered | 0 | 0 
male preterm infant | 0 | 0 
750g | 0 | 0 
neonatal ICU | 0 | 0 
mechanical ventilation | 0 | 0 
gangrenous sigmoid colon | 0 | 0 
ischemic changes | 0 | 0 
necrotic colon | 0 | 0 
posteriorly displaced by pregnant uterus | 0 | 0 
lower segment caesarean section | 0 | 0 
Hartmann’s procedure | 0 | 0 
end colostomy | 0 | 0 
closure of rectal stump | 0 | 0 
post-operative course uneventful | 0 | 216 
discharged home | 216 | 216 
child discharged home | 720 | 720 
reversal of Hartmann’s | 4320 | 4320 
bowel continuity restored | 4320 | 4320 
colo-rectal anastomosis | 4320 | 4320