44 years old | 0
male | 0
admitted to the hospital | 0
weakness | -48
physical deconditioning | -48
type I diabetes mellitus | -6720
peptic ulcer disease | -6720
depression | -6720
seizure disorder | -6720
Charcot foot | -6720
mild developmental delay | -6720
insulin detemir | -6720
escitalopram | -6720
depakote | -6720
clonazepam | -6720
gabapentin | -6720
levetiracetam | -6720
lisinopril | -6720
finasteride | -6720
non-compliance to medications | -6720
history of diabetic ketoacidosis | -6720
substance abuse | -6720
tobacco use | -6720
alcohol use | -6720
marijuana use | -6720
diabetic ketoacidosis | 0
acute kidney injury | 0
acute tubular necrosis | 0
dehydration | 0
hyperkalemia | 0
intravenous fluids | 0
insulin infusion | 0
blood culture | 0
methicillin-susceptible Staphylococcus aureus | 0
vancomycin | 0
piperacillin/tazobactam | 0
persistent positive blood cultures | 24
orthopedic consultation | 24
computerized tomography scan | 24
non-union of left humerus | 8760
osteomyelitis | 24
incision and drainage | 48
drains placed | 48
septicemia | 48
localized abscess | 48
cardiac transthoracic echo | 72
transesophageal echocardiography | 72
benzocaine | 72
lidocaine | 72
hypoxemia | 72
oxygen saturation 85% | 72
arterial blood gas | 72
methemoglobinemia | 72
methylene blue | 72
oxygen saturation 92-94% | 74
repeat methemoglobin levels | 74
hypoxia improved | 74
repeat blood cultures | 96
negative blood cultures | 96
discharged | 120