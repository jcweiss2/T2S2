14 years old | 0
female | 0
obesity | 0
confluent and reticulated papillomatosis | 0
minocycline 100 mg daily | -672
admitted to intensive care unit | 0
acute multiorgan dysfunction | 0
acute kidney injury | 0
hepatic dysfunction | 0
pneumonia | 0
shock | 0
fever | -168
lymphadenopathy | -168
facial edema | -168
minocycline discontinued | -216
broad-spectrum antibiotics administered | -216
condition deteriorated | -168
transferred to academic center | 0
diffuse exanthematous eruption on trunk | 0
pseudovesicular erythematous papules on face, chest, and intertriginous areas | 0
significant facial edema | 0
hyperpigmented, reticulated plaques on chest | 0
Fitzpatrick skin type V-VI | 0
elevated white blood cell (65.0) | 0
eosinophil differential (17%) | 0
elevated creatinine (1.85) | 0
elevated aspartate aminotransferase (2650) | 0
elevated alanine transaminase (767) | 0
elevated alkaline phosphatase (181) | 0
elevated prothrombin time (25.1) | 0
elevated partial thromboplastin time (62.1) | 0
elevated ferritin (9259.2) | 0
elevated lactate dehydrogenase (7326) | 0
elevated procalcitonin (82.18) | 0
elevated fibrin (90) | 0
elevated erythrocyte sedimentation rate (26) | 0
elevated cytokines (IL-2, IL-2R, IL-4, IL-5, IL-6, IL-8, IL-10, IL-13, IL-17, IFN-γ) | 0
elevated human herpesvirus 6 polymerase chain reaction | 0
occult malignancy ruled out | 0
autoimmune and autoinflammatory etiologies evaluated | 0
whole genome sequencing returned negative | 0
human leukocyte antigen testing negative | 0
diagnosed with minocycline-induced DRESS | 0
secondary HLH | 0
RegiSCAR score 7 | 0
high dose steroids (methylprednisolone) | 24
dexamethasone | 72
anakinra | 24
siltuximab | 24
ruxolitinib | 96
total plasma exchange | 72
broad spectrum antibiotics discontinued | 24
recalcitrant hypotension | 0
asystole | 0
passed away | 0
