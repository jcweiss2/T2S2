31 years old | 0
    female | 0
    pancreas-kidney transplant | -87600
    advanced diabetic nephropathy | -87600
    end-stage renal disease | -87600
    chronic renal graft dysfunction | -87600
    regular hemodialysis initiation | -87600
    mycophenolate therapy | 0
    tacrolimus therapy | 0
    prednisolone therapy | 0
    fever | -72
    shortness of breath | -72
    dry cough | -72
    shivering | -72
    high-grade fever | -72
    suspected catheter related blood stream infection | 0
    type 1 diabetes | 0
    hypertension | 0
    bronchial asthma | 0
    glaucoma | 0
    depression | 0
    mild chest discomfort | 0
    temperature 39.4°C | 0
    pulse 112 beats/min | 0
    respiratory rate 24 breaths/min | 0
    oxygen saturation 90% | 0
    blood pressure 138/75 mmHg | 0
    WBC 9.44×10³/μL | 0
    RBC 3.46×10⁶/mcL | 0
    hemoglobin 9.0 g/dL | 0
    neutrophils 86% | 0
    lymphocytes 8% | 0
    absolute neutrophil count 7.17×10³/mcL | 0
    RDW 18.0 | 0
    serum creatinine 541 μmol/L | 0
    urea 11.66 mmol/L | 0
    potassium 4.85 mmol/L | 0
    sodium 139 mmol/L | 0
    phosphorus 2.24 mmol/L | 0
    eGFR 8.4 mL/min/1.73 m² | 0
    total protein 51 g/L | 0
    albumin 23.3 g/L | 0
    CRP 78.0 mg/L | 0
    procalcitonin 3.25 μg/L | 0
    D-dimer 1.40 mg/L | 0
    random blood sugar 7.5 mmol/L | 0
    HbA1C 6.7% | 0
    arterial blood gas pH 7.349 | 0
    pCO2 40.9 mmHg | 0
    pO2 115.4 mmHg | 0
    HCO3 22.0 mmol/L | 0
    chest CT ground glass veiling | 0
    chest CT air space consolidations | 0
    chest CT reticulo-nodular infiltrates | 0
    chest X-ray bilateral multifocal pulmonary opacities | 0
    line related sepsis | 0
    tacrolimus continued | 0
    mycophenolate withheld | 0
    prednisolone increased | 0
    empiric antibiotic therapy | 0
    vancomycin initiated | 0
    meropenem initiated | 0
    amikacin initiated | 0
    regular hemodialysis sessions | 0
    RT-PCR for COVID-19 sent | 0
    blood culture sent | 0
    RT-PCR negative | 24
    blood culture negative | 72
    bronchoscopy refused | 0
    chills | 168
    shivering | 168
    high-grade fever | 168
    desaturating on 15L NRBM | 168
    oxygen saturation 82–83% | 168
    HFNC initiated | 168
    ICU admission | 168
    non-invasive CPAP | 168
    hemodialysis in ICU | 168
    repeat blood cultures sent | 168
    sputum cultures sent | 168
    TB workup sent | 168
    oxygen requirements increased | 168
    chest X-ray bilateral multi-lobar opacities | 168
    hemodialysis in ICU | 168
    alternated between NIV and HFNC | 168
    blood cultures negative | 168
    sputum cultures negative | 168
    TB screen negative | 168
    bronchoscopy refused again | 168
    PCP treatment initiated | 192
    TMP/SMX initiated | 192
    vancomycin stopped | 192
    meropenem stopped | 192
    clinical improvement | 192
    chest X-ray improvement | 192
    sputum PCR positive for Pneumocystis jirovecii | 192
    high-grade fever | 360
    condition deteriorated | 360
    pan-culture sent | 360
    vancomycin restarted | 360
    meropenem restarted | 360
    yeast cells in blood culture | 360
    anidulafungin initiated | 360
    tachypneic | 360
    respiratory rate 40/min | 360
    severe respiratory distress | 360
    chest X-ray bilateral ground glass opacities | 360
    no neurological symptoms | 360
    severe hypoxemia | 360
    unresponsive | 360
    intubation | 360
    mechanical ventilation | 360
    bradycardia | 360
    asystole | 360
    CPR initiated | 360
    death | 360
    blood culture positive for Cryptococcus neoformans | 480
    