51 years old | 0
    male | 0
    Caucasian | 0
    admitted March/April 2009 | 0
    presented with dyspnoea | -672
    presented with abdominal pain | -672
    presented with abdominal distension | -672
    diagnosed with pyelonephritis | -672
    required haemofiltration | -672
    computed tomography scan at diagnosis | -672
    no cardiac changes | -672
    subsequent imaging with CT scan on Day 12 | -576
    cardiomegaly | -576
    moderate-sized pericardial effusion | -576
    diffuse mid-wall myocardial calcification | -576
    transthoracic echocardiogram on Day 32 | -456
    mildly dilated left ventricular | -456
    moderate systolic dysfunction | -456
    pericardial effusion deemed haemodynamically not significant | -456
    LV ejection fraction not quantified | -456
    admitted April 2018 | 0
    presented with cerebrovascular event | -2160
    transthoracic echocardiogram showed severe LV dysfunction | -2160
    LVEF 22% | -2160
    apical thrombus measuring 1.5 cm × 0.9 cm | -2160
    treated with anticoagulation | -2160
    admitted November 2018 | 0
    6-month history of worsening dyspnoea | -4320
    peripheral pitting oedema | -4320
    electrocardiogram showed left atrial enlargement | 0
    electrocardiogram showed inferior pathological Q waves | 0
    transthoracic echocardiogram showed severe LV dysfunction | 0
    LVEF 20% | 0
    commenced on anti-failure medical therapy | 0
    further investigations | 0
    cardiac CT November 2018 | 0
    mild coronary artery disease | 0
    no significant stenosis | 0
    dilated LV | 0
    diffuse LV mid-myocardial calcification | 0
    cardiac magnetic resonance imaging October 2019 | 8760
    diffuse extensive mid-myocardial late gadolinium enhancement | 8760
    moderately dilated LV | 8760
    LVEF 34% | 8760
    continued on anti-failure medical therapy April 2020 | 13560
    stable New York Heart Association class II | 13560
    prophylactic implantable cardioverter-defibrillator implantation | 13560
    presented with worsening dyspnoea over 6 months | 0
    lower leg oedema | 0
    orthopnoea | 0
    paroxysmal nocturnal dyspnoea | 0
    exercise tolerance limited to 40–50 m | 0
    denied chest pain | 0
    denied abdominal pain | 0
    denied palpitations | 0
    denied syncope | 0
    no history of smoking | 0
    no excessive alcohol consumption | 0
    no drug use | 0
    past history of urosepsis nine years prior | -79056
    past history of cerebrovascular event 6 months prior | -4320
    presented with right upper quadrant pain | -79056
    abdominal distension | -79056
    worsening dyspnoea | -79056
    CT scan identified bladder calculus | -79056
    complicated by renal failure | -79056
    required short-term haemofiltration | -79056
    serial blood films showed neutrophilia | -79056
    leucoerythroblastic appearance | -79056
    marked left shift | -79056
    follow-up CT scan April 2009 | -79056
    diffuse LV mid-myocardial calcification | -79056
    transthoracic echocardiogram showed mildly dilated LV | -79056
    no significant pericardial effusion | -79056
    no cardiac symptoms until April 2018 | -2160
    large LV apical thrombus detected | -2160
    bilateral below-knee pitting oedema | 0
    signs of respiratory distress | 0
    heart rate 80 beats/min | 0
    blood pressure 140/90 mmHg | 0
    respiratory rate 18 breaths/minute | 0
    SpO2 98% on room air | 0
    temperature 37.0°C | 0
    not overweight | 0
    no peripheral signs of infective endocarditis | 0
    no respiratory disease | 0
    no hepatic disease | 0
    non-displaced apex beat | 0
    no palpable thrills | 0
    no right ventricular heave | 0
    S1 and S2 heart sounds | 0
    no added sounds | 0
    no murmurs | 0
    no lung crepitations | 0
    ECG showed no acute T wave changes | 0
    ECG showed no acute ST segment changes | 0
    normal cardiac troponin levels | 0
    LVEF quantified at 20% | 0
    serological tests for sarcoidosis normal | 0
    normal serum angiotensin converting enzyme | 0
    normal calcium | 0
    normal phosphate levels | 0
    serological screens for autoimmune pathologies normal | 0
    negative Legionella pneumophila/longbeachae antibodies | 0
    negative Mycoplasma pneumoniae antibodies | 0
    negative Chlamydia antibodies | 0
    negative hepatitis B virus | 0
    negative hepatitis C virus | 0
    negative HIV antibody/antigen combo | 0
    diagnosed with nonAischaemic cardiomyopathy | 0
    commenced on valsartan/sacubitril | 0
    commenced on spironolactone | 0
    commenced on frusemide | 0
    commenced on atorvastatin | 0
    commenced on bisoprolol | 0
    commenced on warfarin | 0
    CMRI October 2019 showed LVEF 34% | 8760
    maintained New York Heart Association class II | 13560
    prophylactic implantable cardioverterAdefibrillator April 2020 | 13560

    