28 years old | 0
male | 0
attended a health center | -24
fatigue | -24
anosmia | -24
dyspnea | -24
SpO2 levels were 55% | -24
nasal cannula oxygen therapy | -24
SpO2 levels improved to 75% | -24
hospitalized | 0
evaluated at an emergency department | 0
chest radiography | 0
bilateral lung infiltrates | 0
RT-PCR swab tested positive for SARS-CoV-2 infection | 0
admitted in a COVID-19 infirmary unit | 0
non-invasive ventilation support | 0
intubation | 0
invasive mechanical ventilation | 0
ventral decubitus positioning | 0
Escherichia coli detected on sputum culture | 48
methicillin-sensitive Staphylococcus aureus detected on sputum culture | 48
superinfection | 48
amoxicillin prescribed | 48
blood culture revealed methicillin-resistant Staphylococcus aureus | 48
methicillin-resistant Staphylococcus aureus dismissed | 48
steady clinical improvement | 72
extubated | 72
discharged | 168
retrosternal thoracalgia | 168
thoracalgia irradiating to the left upper limb | 168
abduction and external rotation limited due to pain | 168
soft tissue swelling of the shoulder and arm | 168
fever | 168
increased levels of C-reactive protein | 168
admitted for further investigation and treatment planning | 168
gentamicin prescribed | 168
gentamicin administered | 168
thoracic CT with intravenous contrast administration | 177
scapulohumeral synovitis | 177
intra-muscular collections | 177
glenohumeral joint fluid | 177
bilateral shoulder magnetic resonance imaging (MRI) with intravenous contrast administration | 180
infraspinatus fossa collections | 180
subscapular fossa collections | 180
capsular thickening | 180
increased signal intensity post-gadolinium administration | 180
septic arthritis | 180
rotator cuff collections | 180
myonecrosis | 180
aspiration of the infraspinatus fossa collection | 192
seropurulent fluid sent for analysis | 192
drainage catheter left on the left infraspinatus collection | 192
drainage catheter removed | 193
improvement of left shoulder range of motion | 216
physical rehabilitation exercises | 216
transferred to another hospital | 216
indication to continue physical therapy and rehabilitation exercises | 216