19 years old | 0
male | 0
Saudi | 0
admitted to the hospital | 0
fever | 0
anaemia | 0
thrombocytopenia | 0
hypercalcemia | 0
normal white cell count | 0
Philadelphia positive ALL | 0
induction chemotherapy | 0
prednisolone | 0
vincristine | 0
idarubicin | 0
Lasparaginase | 0
intrathecal methotrexate | 0
correcting hypercalcemia with intravenous fluids | 0
correcting hypercalcemia with clodronate | 0
fever | -240
diarrhea | -240
E.coli | -240
Klebsiella pneumoniae | -240
intravenous ceftazidime | -240
intravenous amikacin | -240
painful nodule over the left thigh | -504
Pseudomonas aeruginosa | -504
MRSA | -504
E.coli | -504
change ceftazidime and amikacin to imipenem, ciprofloxacin, and vancomycin | -504
central venous catheter removed | -504
induction course of chemotherapy placed on hold | -504
G-CSF initiated | -504
cellulitis | -504
fluid collection | -504
surgical incision and drainage | -504
transferred to the intensive care unit | -504
hemodynamically unstable | -192
ventilatory support | -192
inotropic support | -192
A. xylosoxidans | -192
septic shock | -192
multiorgan failure | -192
intravenous colistin | -192
cardiac arrest | -24
died | 0