34 years old | 0
male | 0
admitted to the hospital | 0
recurrent fever | -3600
rigors | -3600
high fever | -720
chills | -720
right leg pain | -720
lung and soft tissue infections | -720
antibiotics | -720
dyspnea | -718
cough | -718
chest pain | -718
elevation in white blood cell (WBC) counts | -718
high neutrophil percentage | -718
procalcitonin (PCT) level increased | -718
lung infection with encapsulated effusion | -718
abscess in the soft tissues of the right lower leg | -718
incision and drainage of the abscess | -718
antibiotic therapy with ceftazidime | -718
Proteus vulgaris growth | -713
imipenem infusion | -713
sulbactam/cefoperazone infusion | -713
temperature within 37.0 °C | -708
respiratory symptoms improved | -708
leg wound coalesced | -708
recurrent fever | -703
cough | -703
chills | -703
Morganella morganii growth | -696
sulperazone infusion | -696
discharged | -696
fever with chills and cough recurred | -672
antibiotic therapy repeatedly | -672
higher fever | 0
chills | 0
chest pain | 0
cough | 0
fatigue | 0
tachycardia | 0
blood pressure of 108/70 mmHg | 0
temperature of 40.2 °C | 0
respiratory rate of 24 breaths per minute | 0
oxygen saturation of 96% | 0
grade II systolic murmur | 0
normal leukocyte count | 0
elevated neutrophil percentage | 0
CRP level elevated | 0
ESR significantly increased | 0
HIV negative | 0
autoantibodies negative | 0
B lymphocyte count normal | 0
immunoglobulin gamma normal | 0
lymphocyte subpopulations normal | 0
bilateral pulmonary inflammatory shadows | 0
sinus tachycardia | 0
M. morganii growth | 5
NGS confirmed DNA of M. morganii | 5
tricuspid valve vegetation | 5
tricuspid valvuloplasty | 21
vegetation curetted | 21
suspicious perforation not found | 21
bacterial culture of vegetation | 21
M. morganii growth | 21
recovered quickly | 24
pneumonia and fever did not relapse | 96
TTE showed normal heart function | 96
tricuspid valve closed and opened normally | 96
small amount of regurgitation | 96
pulmonary infections completely cured | 120
discharged | 120