52 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
abdominal pain | -48 | 0 | Factual
nausea | -48 | 0 | Factual
vomiting | -48 | 0 | Factual
increased level of liver enzyme alanine aminotransferase | -840 | -840 | Factual
positive autoimmune antibody | -840 | -840 | Factual
elevated immunoglobulin G | -840 | -840 | Factual
coarse liver surface | -840 | -840 | Factual
chronic liver disease | -840 | -840 | Factual
liver biopsy | -840 | -840 | Factual
overlap syndrome | -840 | -840 | Factual
autoimmune hepatitis | -840 | -840 | Factual
ursodeoxycholic acid treatment | -840 | -672 | Factual
prednisolone treatment | -840 | -672 | Factual
reduced prednisolone dose | -672 | -672 | Factual
azathioprine treatment | -672 | 0 | Factual
mild heartburn | -48 | -48 | Factual
abdominal pain worsened | -24 | -24 | Factual
nausea worsened | -24 | -24 | Factual
vomiting worsened | -24 | -24 | Factual
diarrhea | -24 | -24 | Factual
emergency room visit | 0 | 0 | Factual
normal blood pressure | 0 | 0 | Factual
mild fever | 0 | 0 | Factual
tachycardia | 0 | 0 | Factual
tachypnea | 0 | 0 | Factual
abdominal tenderness | 0 | 0 | Factual
reduced white blood cell count | 0 | 0 | Factual
reduced platelet count | 0 | 0 | Factual
decreased neutrophil level | 0 | 0 | Factual
elevated C-reactive protein level | 0 | 0 | Factual
elevated liver enzymes | 0 | 0 | Factual
prothrombin time international normalized ratio | 0 | 0 | Factual
contrast-enhanced abdominal CT | 0 | 0 | Factual
huge stomach with layered wall thickening | 0 | 0 | Factual
air in the stomach wall | 0 | 0 | Factual
decrease of mucosal enhancement | 0 | 0 | Factual
necrotizing gastritis | 0 | 0 | Factual
septic shock | 0 | 0 | Factual
intravenous hydration | 0.5 | 0.5 | Factual
antibiotic treatment | 0.5 | 0.5 | Factual
inotropics | 2 | 2 | Factual
fluid treatment | 2 | 2 | Factual
increased blood pressure | 2 | 2 | Factual
decreased heart rate | 3 | 3 | Factual
stress-induced cardiomyopathy | 3 | 3 | Factual
extracorporeal membrane oxygenation | 3 | 3 | Factual
cardiac arrest | 3 | 3 | Factual
death | 3 | 3 | Factual