18 years old| 0
male | 0
admitted to the hospital | 0
fever | -72
rash | -72
acne |  -672
minocycline |  -672
increased WBC count | 0
eosinophilia| 0
systemic involvement| 0
diffuse erythematous or maculopapular eruption| 0
pruritis | 0
DRESS syndrome | 0
fever persisted | 0
rash persisted | 0
discharged | 24
Separate conjunctive phrases into its component events and assign them the same timestamp (for example, the separation of 'fever and rash' into 2 events: 'fever' and 'rash')  If the event has duration, assign the event time as the start of the time interval. Attempt to use the text span without modifications except 'history of' where applicable. Include all patient events, even if they appear in the discussion; do not omit any events; include termination/discontinuation events; include the pertinent negative findings, like 'no shortness of breath' and 'denies chest pain'.  Show the events and timestamps in rows, each row has two columns: one column for the event, the other column for the timestamp.  The time is a numeric value in hour unit. The two columns are separated by a pipe '|' as a bar-separated file. Skip the title of the table. Reply with the table only. Create a table from the following case:
<|eot_id|><|start_header_id|>user<|end_header_id|>
<|eot_id|><|start_header_id|>assistant<|end_header_id|>
male newborn | 0
transferred to the intensive care unit | 0
respiratory distress | 0
born at 37th gestational week | -24
cesarean section | -24
42-year-old mother | 0
gestational diabetes | -24
poor general appearance | 0
tachycardia | 0
tachypnea | 0
hypotonia | 0
hypoactivity | 0
generalized edema | 0
facial dysmorphic findings | 0
micropenis | 0
tracheal intubation | 0
intratracheal surfactant | 0
severe respiratory acidosis | 0
radiological findings | 0
infant of diabetic mother | 0
respiratory distress syndrome | 0
broad-spectrum antibiotics | 0
umbilical catheterization | 0
peripheral venous puncture prohibited by severe edema | 0
respiratory functions began to improve on third day | 72
continuous positive airway pressure | 72
enteral feeding | 0
no hypoglycemic attack | 0
generalized edema did not diminish | 72
expected weight loss not observed | 72
poor feeding | 72
vomiting | 72
hypoactivity became apparent | 72
hypotonia became apparent | 72
mechanical ventilation again necessary on 7th day | 168
metabolic screening | 168
portal Doppler investigations | 168
splenic Doppler investigations | 168
renal Doppler investigations | 168
echocardiography | 168
central hypothyroidism | 168
low free-thyroxine | 168
slightly elevated thyroid-stimulating hormone | 168
hyponatremia | 168
normal potassium levels | 168
baseline cortisol level 0.44 µg/dL | 168
low-dose adrenocorticotropic hormone test | 168
30th minute cortisol level 4.5 µg/dL | 168
secondary adrenal insufficiency | 168
glucocorticoid replacement with hydrocortisone | 168
thyroid hormone replacement with levothyroxine | 168
vomiting receded | 168
hyponatremia receded | 168
edema significantly improved on third day of treatment | 168
extubated on 15th day | 360
no need for supplemental oxygen on 23rd day | 552
gonadotrophic hormone levels below mini-puberty stage | 552
congenital hypopituitarism | 0
no hypoglycemia | 0
severe respiratory distress | 0
no specific symptom like hypoglycemia | 0
negative acute phase reactants | 0
no response to antimicrobial treatment | 0
slightly elevated TSH | 168
hyponatremia present | 168
baseline cortisol low | 168
no midline alterations | 0
no weight loss | 0
edema diminished | 240
respiratory distress disappeared | 240
enteral feeding | 240
vomiting ceased | 240
hydrocortisone initiated | 168
levothyroxine initiated | 168
ampicillin+gentamicin | 0
vancomysin+meropenem | 168
extubation | 360
no supplemental oxygen needed | 552
<|begin_of_text|>
<|start_header_id|>system<|end_header_id|>
