50 years old | 0
male | 0
admitted to the hospital | 0
dry cough | -96
chills | -96
fever | -96
back pain | -96
cough | -96
visited another clinic | -96
prescribed acetaminophen | -96
prescribed carbocysteine | -96
no gastrointestinal symptoms | -96
no diarrhea | -96
20-pack-year smoker | 0
does not drink alcohol | 0
lives in an over 40-year-old house | 0
contaminated shower use presumed | 0
works in a bar | 0
does not use a humidifier or an air conditioner | 0
no recent history of travel to a spa or other countries | 0
on maintenance HD for three years | 0
diabetic kidney disease | 0
percutaneous coronary intervention of his right coronary artery | -2880
angina pectoris | -2880
congestive heart failure | 0
taking beta blockers | 0
taking angiotensin receptor blockers | 0
echocardiography showed an ejection fraction of 33% | -672
diffuse hypokinesis | -672
echocardiography on admission revealed an ejection fraction of 30% | 0
no history of gastrointestinal disorders | 0
no family history of diabetes | 0
no family history of HD | 0
no family history of immunodeficiency | 0
body temperature of 38.9 °C | 0
blood pressure of 131/97 mmHg | 0
heart rate of 117 per minute | 0
respiratory rate of 18 per minute | 0
arterial oxygen saturation on pulse oximetry was 96% | 0
consciousness was intact | 0
left pulmonary rales | 0
bilateral lower leg edema | 0
no xerostomia | 0
elevated leukocyte count | 0
markedly elevated C-reactive protein levels | 0
severe abnormalities in the liver function | 0
severe abnormalities in creatine kinase value | 0
moderate hypoxemia | 0
tachycardia | 0
no specific ST elevation to indicate ischemic heart disease | 0
lobular infiltrates in the left lower lung field | 0
mild heart enlargement | 0
no significant amount of pleural effusion | 0
lobar consolidation with areas of air bronchogram in the left lower lobe | 0
chronic liver injury | 0
fatty liver | 0
bacterial pneumonia with severe liver dysfunction diagnosed | 0
A-DROP score <1 | 0
quick Sequential Organ Failure Assessment score 0 | 0
started piperacillin/tazobactam | 0
lab results worsened | 24
started oral azithromycin | 24
consciousness level and systolic blood pressure deteriorated | 34
diagnosed with septic shock | 34
started intravenous infusion of noradrenaline | 34
developed bradycardia | 48
cardiac arrest | 48
started cardiopulmonary resuscitation | 48
defibrillation attempts | 48
adrenaline bolus doses | 48
transferred to the intensive-care unit | 48
started hydrocortisone phosphate | 48
started gamma globulin | 48
started continuous renal replacement therapy | 72
reduced noradrenaline dose | 72
changed oral azithromycin to levofloxacin | 72
blood pressure suddenly dropped | 120
discontinued CRRT | 120
died | 120
Legionella pneumophila serotype 1 detected on sputum multiplex PCR | 120
autopsy showed lobar pneumonia | 120
hepatic lobular central congestion and shock liver | 120
yellow pleural effusion | 120
no pleural adhesion | 120
centrilobular congestion and necrosis without an inflammatory response | 120
no new heart infarctions | 120
afferent cardiac hypertrophy due to hypertension | 120
lower limb ischemia | 120