5 weeks old | 0
infant | 0
male | 0
admitted to the Emergency Room | 0
fever | 0
fussiness | 0
born at 40 weeks gestation | -672
C-section | -672
failure to progress | -672
G1P1 mother | -672
negative prenatal serologies | -672
APGAR scores were 8 and 9 | -672
hypoglycemia | -672
respiratory distress | -672
tachypnea | -672
resolved by day 2 of life | -48
newborn screening test was positive for congenital adrenal hyperplasia | -48
Pediatric endocrinology was consulted | -48
cortisol level obtained on day 2 of life was 1.2 mcg/dL | -48
17-hydroxyprogesterone was 813 ng/dL | -48
ACTH stimulation test was performed | -48
17 hydroxyprogesterone level of 17 836 ng/dl | -48
cortisol level of 3.9 mcg/dl | -48
initiated on hydrocortisone therapy | -48
fludrocortisone 0.1 mg daily | -48
Sodium chloride 2 grams divided in several feedings | -48
father reported symptoms of cough and a runny nose | -24
presented to the ER with fever and increased fussiness | 0
no respiratory distress | 0
no diarrhea | 0
no vomiting | 0
no rash | 0
no decreased feeding | 0
afebrile | 0
oxygen saturation of 100% | 0
irritable | 0
skin was mottled | 0
no chest retractions | 0
no tachypnea | 0
no nasal flaring | 0
WBC 7.2 bil/L | 0
neutrophils 2.1 bil/L | 0
lymphocytes 2.5 bil/L | 0
monocytes 2 bil/L | 0
Na 136 mmol/L | 0
potassium 5.9 mmol/L | 0
HCO3 22 mmol/L | 0
glucose of 110 mg/dL | 0
BUN 8 mg/dL | 0
creatinine 0.33 mg/dL | 0
CRP 1.9 mg/L | 0
SARS-CoV-2 by Nucleic Acid Amplification was detected | 0
blood culture was negative | 0
urinalysis was negative | 0
urine culture was negative | 0
chest x-ray demonstrated mild streaky bilateral perihilar streaks | 0
placed on triple maintenance hydrocortisone | 0
fludrocortisone 0.15 mg daily | 0
received a normal saline bolus | 0
placed on maintenance IV fluids | 0
transferred to the Pediatric Intensive Care Unit | 0
Pediatric infectious disease specialists were consulted | 0
remained hemodynamically stable | 24
fed appropriately | 24
did not require respiratory support | 24
discharged | 48
stress hydrocortisone dose was weaned down | 48
doing well | 336