72 years old | 0
male | 0
cirrhosis | 0
hepatocellular carcinoma | 0
systemic immunotherapy | 0
tocilizumab | 0
atezolizumab | 0
bevacizumab | 0
oral prednisone | 0
systemic inflammatory response | 0
presented to the emergency department | -312
confusion | -312
lethargy | -312
bilateral lower extremity edema | -312
recurrent falls | -312
lacerations | -336
dog lick | -336
hospital admission | 0
feeling unwell | 0
described as being in bad shape | 0
temperature of 100.0°F | 0
blood pressure of 85/50 | 0
heart rate in the 80s | 0
increasing confusion | 0
red leg ulceration | 0
hot leg ulceration | 0
painful leg ulceration | 0
elevated white blood cell count | 0
left shift | 0
sepsis protocol initiated | 0
admitted to the intensive care unit | 0
broad-spectrum antimicrobials initiated | 0
vancomycin | 0
piperacillin/tazobactam | 0
acute kidney injury | 24
antimicrobials changed to vancomycin | 24
cefepime | 24
metronidazole | 24
bacterial culture specimens obtained | 0
blood cultures drawn | 0
cultures positive for M. canis | 24
Staphylococcus aureus | 24
clinical improvement observed | 72
repeat blood cultures negative | 72
fever resolved | 72
leg wounds improved | 72
white blood cell count trended downwards | 72
neutrophil counts trended downwards | 72
IV cefepime continued for five days | 72
oral cefdinir | 312
outpatient therapy | 312
