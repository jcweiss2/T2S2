68 years old|0
male|0
diabetes mellitus type II|0
hypertension|0
chronic kidney disease stage 5|0
heart failure with preserved ejection fraction (Grade III)|0
admitted to the hospital|0
shortness of breath|0
generalized body aches|0
worsening kidney function|0
serum creatinine 245 umol/L|-720
hemodialysis|264
hypotension 87/57 mmHg|528
lethargic|528
decreased urine output|528
shifted to MICU|528
crystalloids bolus|528
norepinephrine infusion|528
echo on day 22|528
moderate pericardial effusion|528
increased risk of bleeding|528
INR 1.7|528
FFP 4 units|528
increased vasopressors requirements|552
lactate 8 mmol/L|552
anuric|552
continuous renal replacement therapy|552
increased ALT to 1729 U/L|552
increased AST to 1772 U/L|552
INR 2|552
acute ischemic hepatitis|552
coagulopathy|552
emergency pericardiocentesis|552
FFP 4 units|552
vitamin K 10 mg|552
cardiac index 0.9 L/min/m2|552
systemic vascular resistance >4000 dynes/sec/cm5|552
cardiogenic shock|552
cardiac tamponade|552
INR 2.3|552
FEIBA 2500 units|552
INR 1.9|552
pericardiocentesis|552
draining 60 mL fluid|552
hemodynamic deterioration|624
asystole cardiac arrest|624
cardiopulmonary resuscitation|624
death|624
