66 years old | 0  
    woman | 0  
    advanced diffuse large B-cell lymphoma (DLBCL) | 0  
    referred for CAR T cell therapy | 0  
    diagnosed with DLBCL | -52560  
    no significant past medical history | -52560  
    received 10 cycles of R-CHOP | -52560  
    lifetime exposure of doxorubicin >500 mg/m2 | -52560  
    autologous hematopoietic stem cell transplant | -52560  
    DLBCL recurred | -35040  
    6 more cycles of R-CHOP | -35040  
    transthoracic echocardiogram (TTE) | -720  
    LVEF 55% to 60% | -720  
    global longitudinal strain −12% | -720  
    admitted to the hospital | 0  
    acute decompensated heart failure (HF) | 0  
    repeat TTE | 0  
    LVEF 25% | 0  
    global left ventricular (LV) dysfunction | 0  
    positron emission tomography scan imaging demonstrated progression of DLBCL | 0  
    new pulmonary nodules | 0  
    referred to our center for consideration of CAR T cell therapy | 0  
    coronary computed tomography demonstrated mild coronary artery disease | 0  
    cardiac magnetic resonance imaging showed no evidence of infiltrative or inflammatory disease | 0  
    presumed to have anthracycline-induced cardiomyopathy | 0  
    initiated on furosemide | 0  
    initiated on GDMT | 0  
    lisinopril 2.5 mg | 0  
    metoprolol succinate 12.5 mg daily | 0  
    up-titration of GDMT limited | 0  
    spironolactone or eplerenone could not be added | 0  
    hypotension | 0  
    referred to cardio-oncologist for risk stratification prior to CAR T cell therapy | 0  
    good exercise tolerance | 0  
    riding stationary bike | 0  
    right heart catheterization (RHC) | 0  
    mildly elevated biventricular filling pressures | 0  
    normal cardiac output | 0  
    right atrium 10 mm Hg | 0  
    pulmonary artery 36/20/27 mm Hg | 0  
    pulmonary capillary wedge pressure 16 mm Hg | 0  
    Fick cardiac output 5.1 l/min | 0  
    Fick cardiac index 2.9 l/min/m2 | 0  
    mixed venous oxygen saturation 57.4% | 0  
    multidisciplinary discussions held | 0  
    decision for 3-month trial of GDMT | 0  
    concern for CRS during CAR T cell therapy | 0  
    manifestations of CRS | 0  
    fevers | 0  
    derangements in blood pressure | 0  
    derangements in oxygenation | 0  
    hypotension | 0  
    hypoxemia | 0  
    vasodilatory shock requiring vasopressors | 0  
    severe hypoxemia necessitating intubation | 0  
    hypoxemia from capillary leak syndrome | 0  
    low-pressure pulmonary edema | 0  
    atrial arrhythmias | 0  
    ventricular arrhythmias | 0  
    ventricular dysfunction | 0  
    invasive pulmonary artery catheter monitoring considered | 0  
    risk of infection prohibitive | 0  
    lympho-depleting chemotherapy prior to CAR T cell therapy | 0  
    decision to implant CardioMEMS device | 0  
    after 3 months of GDMT | 720  
    repeat RHC | 720  
    normal filling pressures | 720  
    preserved cardiac output | 720  
    right atrium 2 mm Hg | 720  
    pulmonary artery 25/12/18 mm Hg | 720  
    pulmonary capillary wedge pressure 15 mm Hg | 720  
    Fick cardiac output 4.7 l/min | 720  
    Fick cardiac index 2.8 l/min/m2 | 720  
    mixed venous oxygen saturation 61.5% | 720  
    placement of CardioMEMS device | 720  
    repeat TTE | 720  
    LVEF 24.6% | 720  
    right ventricular performance improved | 720  
    admitted for pre-treatment with lympho-depleting chemotherapy | 792  
    fludarabine | 792  
    cyclophosphamide | 792  
    neutropenic fever | 792  
    hypotension | 792  
    started on intravenous antibiotics | 792  
    GDMT held | 792  
    infusion of axicabtagene ciloleucel CAR T cells | 816  
    developed mild CRS | 864  
    fevers | 864  
    sinus tachycardia to 150s | 864  
    systolic blood pressures in 90s | 864  
    CardioMEMS demonstrated PAd 20 mm Hg | 864  
    given intravenous furosemide 20 mg | 864  
    given tocilizumab | 864  
    day 3 | 864  
    worsening tachypnea | 864  
    new oxygen requirement | 864  
    second dose of tocilizumab | 864  
    chest x-ray diffuse pulmonary opacities | 864  
    PAd 10 mm Hg | 864  
    noncardiogenic pulmonary edema | 864  
    held diuretic agents | 864  
    monitoring volume status | 864  
    oncology nurses performed CardioMEMS measurements | 864  
    advanced HF consult service rounded daily | 864  
    day 6 | 960  
    atrial flutter | 960  
    rapid ventricular rates | 960  
    acute hypoxic respiratory failure | 960  
    cardiogenic pulmonary edema | 960  
    PAd 23 mm Hg | 960  
    required intubation | 960  
    initiated on low-dose norepinephrine | 960  
    started on amiodarone | 960  
    converted to sinus rhythm | 960  
    intermittent doses of intravenous furosemide 20 to 40 mg | 960  
    PAd between 10 to 20 mm Hg | 960  
    weaned off vasopressors | 960  
    extubated | 960  
    daily discussions | 960  
    completed CAR T cell therapy | 1440  
    discharged to acute rehabilitation | 1440  
    one-month hospitalization | 1440  
    unable to restart GDMT | 1440  
    hypotension | 1440  
    PAd 6 mm Hg at discharge | 1440  
    plan for positron emission tomography scan | 1440  
    initial course at facility uncomplicated | 1440  
    participated in physical therapy | 1440  
    weekly appointments in oncology clinic | 1440  
    appointment with advanced HF team | 1440  
    rehabilitation providers transmitted CardioMEMS readings | 1440  
    furosemide 20 mg daily restarted | 1440  
    PAd 18 mm Hg | 1440  
    physician reported doing well | 1440  
    15 days later | 1560  
    acute shortness of breath | 1560  
    oxygen saturation 88% | 1560  
    no dyspnea prior | 1560  
    nausea for past 3 days | 1560  
    taken by ambulance | 1560  
    chest x-ray pulmonary edema | 1560  
    possible left lower lobe infiltrate | 1560  
    PAd 22 mm Hg | 1560  
    intubated | 1560  
    progressive hypoxic respiratory failure | 1560  
    bedside TTE showed severe LV dysfunction | 1560  
    normal right ventricular function | 1560  
    treated with multiple vasopressors | 1560  
    mixed septic and cardiogenic shock | 1560  
    cardiac arrest | 1560  
    ventricular tachycardia | 1560  
    expired | 1560  
    