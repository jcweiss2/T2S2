58 years old | 0
female | 0
internal haemorrhoids | 0
undergoes rubber-band ligation (RBL) | 0
osteoporosis | 0
dyslipidemia | 0
depression | 0
pelvic pain | 48
dysuria | 48
no necrosis | 48
no signs of infection | 48
empirical intravenous antibiotics | 48
ciprofloxacin | 48
metronidazole | 48
clinical observation | 48
condition did not improve | 48
white blood count (WBC) increased significantly (24,000/μL) | 48
transferred to a referral centre | 48
band removed | 48
small superficial abscess drained | 48
computed tomography (CT) scan of the abdomen and pelvis | 48
rectosigmoiditis | 48
moderate to severe amount of ascites | 48
no pneumatosis | 48
exploratory laparoscopy performed | 48
important amount of serous ascites | 48
severe systemic inflammatory response syndrome (SIRS) | 48
required intensive care | 48
clinical deterioration | 48
persistent leukocytosis (25,000/μL) | 48
transferred to tertiary care centre | 48
suspicion of ischaemic colitis | 48
hemodynamic deterioration | 48
respiratory deterioration | 48
ventilator support | 48
acute respiratory distress syndrome (ARDS) | 48
antibiotics’ spectrum broadened to carbapenem | 48
colonoscopy to mid-transverse colon performed | 48
superficially necrotic 2 cm segment in lower rectum | 48
petechial mucosa | 48
inotropic support with vasopressors | 72
aggressive volemic resuscitation | 72
ventilator support | 72
antibiotics | 72
modest improvement | 72
WBC count decreased from 30,000 to 23,000/μL | 72
repeat abdominopelvic CT scan | 96
circumferential thickening of rectosigmoid colon | 96
no pneumatosis | 96
state of shock subsided | 96
extubated | 216
transferred to floor | 216
discharged from hospital | 216
recovered from intensive care unit myopathy | 216
recovered from prolonged intubation | 216
intensive rehabilitation | 216
muscular weakness | several months
poor exercise tolerance | several months
colonoscopy performed (follow-up) | 26280
normal colonoscopy | 26280
followed by respirologist | 26280
persistent dyspnea | 26280
improving dyspnea | 26280
severe deconditioning during hospital stay | 26280
no residual cardiorespiratory injury | 26280
three years after events | 26280
pelvic sepsis | 0
shock | 0
multiple organ failure (MOF) | 0
