21 years old | 0
female | 0
Caucasian | 0
admitted to the obstetric department | 0
pre-term labor | 0
received 10 mg of nifedipine 4 times in 1 hour | 0
pulmonary edema | 0
hypoxemia | 0
transfer to the intensive care unit | 0
blood pressure 101/61 mm Hg | 0
ECG revealed sinus tachycardia (142 bpm) | 0
oxygen saturation 98% under 100% high flow oxygenation | 0
loud first heart sound | 0
diastolic murmur | 0
bilateral wheezing | 0
jugular venous distension | 0
fall in systolic blood pressure | 0
worsening desaturation (78%) | 0
metabolic acidosis | 0
hyperlactatemia (34 mg/dL) | 0
intubated | 0
ventilated (volume-controlled ventilation with FiO2 100% and PEEP at 15 cm H2O) | 0
chest X-ray confirmed pulmonary edema | 0
cardiac echography revealed severe mitral stenosis | 0
normal left ventricular function | 0
enlargement of the left atrium | 0
pressure overload of the left atrium | 0
severe pulmonary hypertension (estimated PAP = 85 mm Hg) | 0
diagnosis of cardiogenic shock precipitated by nifedipine | 0
unknown severe mitral stenosis | 0
administered loop diuretics (furosemide) | 0
administered full-dose heparin | 0
blood pressure stabilized | 0
ultrasound examination showed no fetal distress | 0
transoesophageal echocardiography showed severe rheumatic mitral stenosis (valve area 0.5 cm2, mean gradient 25 mmHg) | 0
Wilkins score 8 | 0
authorization of percutaneous valvuloplasty | 0
spontaneous vaginal delivery | 0
baby alive | 0
transfer to intensive neonatal care unit | 0
mother in critical state with hypotension | 0
needed ventilation | 0
delivery complicated by endometritis | 0
sepsis | 0
treated with ceftriaxone | 0
treated with ampicillin | 0
valvuloplasty postponed | 0
resolution of the infection | 168
percutaneous double balloon mitral valvuloplasty performed | 168
mitral mean gradient reduced from 10 to 3 mmHg | 168
mitral area increased from 0.5 to 1.65 cm2 | 168
pulmonary pressure normalized | 168
rapid recovery | 192
extubated | 192
