18 years old| 0
male| 0
admitted to the hospital| 0
acute respiratory failure due to COVID-19 pneumonia| 0
mechanical ventilation support| 0
mortality rate high| 0
early prone position application| 0
neuromuscular blockers| 0
low tidal volume administration| 0
improved PaO2/FiO2 ratio| 0
decreased mortality| 0
awake prone position combined with noninvasive mechanical ventilation| 0
nasal high-flow applications| 0
corrected ventilation/perfusion incompatibility| 0
provided lung drainage| 0
study conducted| 0
local ethics committee approval| 0
Ministry of Health approval| 0
Clinical Trials registration| 0
informed consent obtained| 0
patients >18 years old included| 0
conventional oxygen therapy with nonrebreather mask oxygen| 0
excluded patients with invasive mechanical ventilation| 0
respiratory acidosis (pH <7.30 and PaCO2 >50 mmHg)| 0
PaO2/FiO2 ratio <150| 0
Glasgow Coma Scale score <12| 0
hemodynamic instability| 0
excluded primary pulmonary pathologies (lung cancer, cardiopulmonary edema, Kartagener’s syndrome)| 0
excluded nasal high-flow therapy| 0
excluded awake PP <12 hours/day| 0
COVID-19 diagnosed with polymerase chain reaction test| 0
pneumonia diagnosed with clinical results and computed tomography findings| 0
acute respiratory failure defined as PaO2/FiO2 ratio <300| 0
FiO2 calculation used| 0
APP group (awake PP 12–18 hours/day)| 0
non,APP group (no awake PP)| 0
recorded demographic data and comorbidities| 0
SpO2, PaO2/FiO2, pH, PaCO2, PaO2 recorded| 0
conventional oxygen therapy administered| 0
SpO2 >93% targeted| 0
awake PP applied intermittently 12–18 hours/day| 0
treatment failure defined as PaO2/FiO2 <150, SpO2 <93%, Glasgow Coma Scale <12, respiratory acidosis| 0
intubation and invasive mechanical ventilation on treatment failure| 0
intubation need recorded| 0
ventilator-free days recorded| 0
ICU stay length recorded| 0
short-term mortality recorded| 0
statistical analysis performed| 0
225 patients examined| 0
61 patients already intubated excluded| 0
36 patients excluded due to respiratory acidosis, low PaO2/FiO2, low Glasgow Coma Scale, hemodynamic instability| 0
52 patients excluded due to nasal high-flow therapy| 0
24 patients excluded due to <12 hours/day awake PP| 0
4 patients excluded due to lung cancer| 0
48 patients included| 0
APP group: 25 patients| 0
non,APP group: 23 patients| 0
APP group lower median age| 0
no significant difference in sex, BMI, comorbidities| 0
initial SpO2, pH, PaO2, PaO2/FiO2 similar| 0
higher initial PaCO2 in APP group| -24
24th hour higher SpO2 and PaO2 in APP group| 24
no significant difference in pH, PaCO2, PaO2/FiO2 at 24th hour| 24
SpO2 increase in APP group| 24
PaO2 increase in APP group| 24
PaCO2 decrease in APP group| 24
pH decrease in non,APP group| 24
ventilator-free days higher in APP group| 24
ICU stay similar| 24
lower intubation requirement in APP group| 24
lower short-term mortality in APP group| 24
acute respiratory failure prevalence ~19%| 0
oxygen treatment requirement 14%| 0
ICU admission risk factors: age >60, male, diabetes, immunodeficiency| 0
mortality risk factors: cardiovascular disease, chronic respiratory disease, diabetes| 0
ARDS assessment| 0
L and H phenotypes identified| 0
PP recommended >12 hours/day| 0
Surviving Sepsis Campaign recommends PP 12–16 hours| 0
PP application difficulties in intubated patients| 0
awake PP preferred in COVID-19| 0
Caputo et al. study: 50 patients, PP improved SpO2| 0
intubation requirement 24%| 0
case report: awake PP with nasal high flow improved PaO2/FiO2| 0
self-PP success in Jiangsu Province| 0
mortality rate 30–40% in ICU, 90% with invasive ventilation| 0
study limitations: not prospective randomized| 0
conclusion: awake PP improves oxygenation, reduces intubation and mortality| 0
no conflicts of interest declared| 0
