30 years old | 0
female | 0
bilateral liposuction | -10
unbearable pain | -10
erythema | -10
blisters | -10
admitted to hospital | 0
febrile | 0
heart rate 128 beats/minute | 0
swelling | 0
tenderness | 0
sutures removed | 0
urine black | 0
leukocytosis | 0
elevated C-reactive protein | 0
elevated serum creatinine | 0
elevated blood urea nitrogen | 0
fasciotomy | 0
drainage | 0
vancomycin | 0
meropenem | 0
sepsis | 0
renal insufficiency | 0
shock | 0
transferred to surgical intensive care unit | 0
continuous renal replacement therapy | 0
anti-infection treatment | 0
blood transfusion | 0
shock correction | 0
exudation | 24
local swelling | 24
extensive fasciotomy | 24
osteofascial compartment incision | 24
vacuum sealing drainage | 24
degeneration | 24
necrosis | 24
high-sensitivity troponin elevated | 24
bilateral iliolumbar local skin edema | 120
inflammatory reaction | 120
subcutaneous effusion | 120
thigh necrotizing fasciitis incision | 120
dilatation | 120
VSD | 120
Candida dubliniensis detected | 120
Klebsiella pneumoniae detected | 120
skin necrotizing area stable | 168
debridement | 168
necrosis | 168
local tissue lacked elasticity | 168
VSD | 168
wounds stable | 168
granulation tissue growth | 168
debridement and skin grafting | 216
skin grafts survived | 216
function of lower limbs recovered | 216
systemic MODS | 0
multiple operations | 0
active treatment | 0
plastic surgery | 0
organ function recovered | 216
discharged | 360