13 years old | 0  
    girl | 0  
    DiGeorge syndrome | 0  
    neonatal truncus arteriosus repair | -109248 (approx. 13 years before admission)  
    severe left pulmonary artery hypoplasia | 0  
    methicillin-sensitive staphylococcal bacteremia | -72 (assuming presentation a few days before admission)  
    infective endocarditis | -72  
    septic pulmonary emboli | -72  
    bilateral pyelonephritis | -72  
    septic shock | -72  
    worsening respiratory failure | -72  
    pulmonary hemorrhage | -72  
    placed on venovenous extracorporeal membrane oxygenation | -72  
    acute hemorrhage around and in the right chest tube | -168 (6 days after ECMO placement, assuming ECMO started at -72, so -72 + 6*24 = 72, but since events before admission, likely timestamp -168)  
    acute hemorrhage in the endotracheal tube | -168  
    computed tomography angiography | -168  
    patent conduit between the right ventricle and the pulmonary artery | 0  
    acute right hemothorax | -168  
    19-mm bilobed presumed mycotic aneurysm | -168  
    extravasation from an intercostal artery | -168  
    placed under general anesthesia | 0  
    perfusionist team support for ECMO | 0  
    left common femoral vein access | 0  
    micropuncture set used | 0  
    9-French Flexor sheath placement | 0  
    7-French APC catheter used | 0  
    digital subtraction arteriography | 0  
    patent pulmonary artery conduit | 0  
    19-mm bilobed mycotic aneurysm confirmed | 0  
    guiding sheath advanced into right pulmonary artery | 0  
    5-French vertebral tip catheter used | 0  
    angled tip Glidewire used | 0  
    cannulation of branch vessel feeding aneurysm | 0  
    decision to occlude aneurysm using balloon occlusion technique | 0  
    Scepter C Occlusion Balloon Catheter placement | 0  
    Synchro 0.014-inch wire used | 0  
    occlusion balloon inflated to 5 mm | 0  
    dead space primed with dimethyl sulfoxide | 0  
    EVOH (Onyx 34) injection | 0  
    mycotic aneurysm filled completely | 0  
    balloon deflated | 0  
    repeat pulmonary arteriography | 0  
    occlusion of mycotic aneurysm | 0  
    preserved flow to normal lung parenchyma | 0  
    right femoral arterial access | 0  
    thoracic aortogram | 0  
    extravasation from right intercostal artery | 0  
    intercostal artery treated with coils and Gelfoam | 0  
    total procedure time 132 minutes | 0  
    returned to pediatric intensive care unit | 0  
    hemorrhage resolved in right chest tube | 24  
    hemorrhage resolved in endotracheal tube | 24  
    care withdrawn due to neurologic deterioration | 96 (3 days after procedure)  
    family declined autopsy | 96  

<|eot_id|>
