73 years old | 0
male | 0
South Asian ethnicity | 0
admitted to the hospital | 0
prior diagnosis of progressive chronic kidney disease | -1300
obstructive uropathy | -1300
recurrent urosepsis | -1300
hydronephrotic left kidney | -1300
insertion of a J-J ureteric stent | -1300
type 2 diabetes mellitus | -1300
ischaemic heart disease | -1300
myocardial infarction | -1300
hypertension | -1300
no history of cardiac dysrhythmia | 0
no prothrombotic diathesis | 0
no cerebrovascular disease | 0
no family history of renal or cerebrovascular disease | 0
not on maintenance antiplatelet agents | 0
not on oral anticoagulants | 0
non-smoker | 0
does not consume alcohol | 0
emergency admission to the intensive care unit | -78
pulmonary oedema | -78
oliguria | -78
serum creatinine of 10.2 mg/dL | -78
established on maintenance thrice weekly HD | -78
right internal jugular tunnelled cuffed central venous catheter | -78
presentation with acute stroke | 0
acute right hemiparesis | 0
aphasia | 0
duration of symptoms 90-min | 0
routine HD 24-h prior to presentation | -24
no complications prior to presentation | -24
blood pressure 190/87 mmHg | 0
capillary blood glucose 86.5 mg/dL | 0
Glasgow Coma Score 15/15 | 0
sinus rhythm on electrocardiogram | 0
urgent CT scan of brain | 0
acute ischaemic stroke | 0
superior parasagittal cortex of the left frontal lobe | 0
no evidence of intracranial haemorrhage | 0
transferred to acute stroke centre | 0
blood pressure 176/75 mmHg | 0
mild right facial droop | 0
right hemiparesis | 0
increased muscle tone in upper limb | 0
lower limb hyper-reflexia | 0
upgoing plantar response in lower limb | 0
dysphasic with receptive and expressive elements | 0
no cardiac murmurs or carotid bruits | 0
clinically euvolaemic | 0
calculated total NIH stroke score 8 | 0
laboratory examinations | 0
Haemoglobin 15.9 g/dL | 0
Total leucocyte count 7.5 × 10^9/mL | 0
Platelet count 161 × 10^9/mL | 0
Sodium 136 mmol/L | 0
Potassium 4.7 mmol/L | 0
Urea 12.2 mmol/L | 0
Creatinine 462 μmol/L | 0
Albumin 44 g/L | 0
Total cholesterol 2.2 mmol/L | 0
C-reactive protein 2 mg/L | 0
INR 1.1 | 0
APTT 27.8 s | 0
Fibrinogen 4.00 g/L | 0
no absolute contraindications to thrombolysis | 0
eligible for trial enrolment | 0
informed consent | 0
randomization | 0
received 54 mg rtPA | 4
rtPA delivery | 4
repeat CT brain scan | 28
small area of haemorrhagic transformation | 28
no other interval change | 28
clinically stable | 28
required sodium valproate | 28
required clobazam | 28
intermittent left upper limb myoclonus | 28
echocardiography | 28
borderline left ventricular hypertrophy | 28
24-h Holter | 28
sinus rhythm with a 1-h paroxysm of asymptomatic atrial fibrillation | 28
no significant carotid stenosis | 28
transferred to specialist renal stroke rehabilitation unit | 96
inpatient for a month | 96
power in upper limb improved | 672
power in lower limb improved | 672
dysphasia improved | 672
residual mild expressive deficit | 672
discharged home | 672
maintenance HD | 672