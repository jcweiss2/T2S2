72 years old | 0
    male | 0
    type-2 diabetes | 0
    diabetic microvascular complications | 0
    diabetic macrovascular complications | 0
    presented with 3-day history of painful left lower leg | -72
    red left lower leg | -72
    swollen left lower leg | -72
    hyperthermic left lower leg | -72
    Co-Amoxicillin commenced by GP | -72
    hospitalized at regional general hospital | 0
    hemodynamically stable | 0
    left foot badly swollen | 0
    left lower leg badly swollen | 0
    tender left foot | 0
    tender left lower leg | 0
    macerated skin in interdigital spaces | 0
    fissures in interdigital spaces | 0
    foot pulses not palpable | 0
    ankle brachial index 0.8 bilaterally | 0
    mild arterial perfusion deficit | 0
    pallanaesthesia | 0
    reduced monofilament sensation | 0
    impaired nociception | 0
    ear-temperature 37.6°C | 0
    BP 161/86 mmHg | 0
    pulse 96/min | 0
    CRP 182 mg/L | 0
    leukocytes 15.2 g/L | 0
    86% neutrophils | 0
    eGFR 80 mL/min/1.73 m2 | 0
    HbA1c 90 mmol/mol | 0
    x-ray showed normal osseous structures | 0
    minimal effusion in left upper ankle joint | 0
    MRI showed bone marrow edema | 0
    bone marrow edema in ankle joint | 0
    bone marrow edema in tarsus | 0
    bone marrow edema in metatarsus | 0
    skin biopsy performed | 0
    histological diagnosis of stasis dermatitis | 0
    antibiotic therapy changed to Amoxicillin/clavulanic acid | 0
    antibiotic therapy changed to Piperacillin/Tazobactam | 0
    discharged | 0
    presented in January 2019 with acute pain in both distal legs | 72
    electrifying pain in left medial malleolus | 72
    bilateral lower extremity edema | 72
    inflammatory signs on left lower leg | 72
    afebrile | 72
    hemodynamically stable | 72
    CRP 28 mg/L | 72
    leukocytes within normal limits | 72
    cellulitis diagnosed | 72
    Co-Amoxicillin started | 72
    painless second-degree ulcer on right fifth MTP joint | 72
    clinical examination | 72
    pulmonary x-ray | 72
    BNP 1341 ng/L | 72
    cardiac decompensation | 72
    treated with diuretics | 72
    x-ray ruled out osteomyelitis of right foot | 72
    MRI ruled out osteomyelitis of right foot | 72
    calcified pedal arteries on x-ray | 72
    mediastinal sclerosis | 72
    vascular review ordered | 72
    reduced toe pressures | 72
    pathologic pulse wave forms | 72
    compromised arterial blood flow | 72
    angiography performed | 72
    percutaneous transluminal angioplasty performed | 72
    discharged after 14 days | 72
    referred to diabetic foot clinic | 72
    wound management | 72
    offloading of right MTP fifth joint | 72
    lesion lateral to right MTP fifth joint | 72
    no adequate progress | 72
    severe pain in left foot | 72
    mild erythema on left foot | 72
    moderate swelling on left foot | 72
    hyperthermia on left foot | 72
    progressive deformity of left ankle joint | 72
    ulcerous lesion with purulent drainage over left lateral malleolus | 72
    large wound cavity probed to bone | 72
    x-ray confirmed complete destruction of left upper ankle joint | 72
    dislocation of left upper ankle joint | 72
    vital signs: auricular temperature 37.8°C | 72
    BP 111/59 mmHg | 72
    pulse rate 74/min | 72
    CRP 68 mg/L | 72
    leukocytes 6.9 G/L | 72
    81.5% neutrophils | 72
    eGFR 40 mL/min/1.73 m2 | 72
    hospitalized | 72
    complete bed rest | 72
    antibiotic therapy with Co-Amoxicillin | 72
    blood cultures showed staphylococcus aureus bacteraemia | 72
    antibiotic regimen changed to Cefazolin | 72
    acute kidney injury | 72
    hemodynamic dysfunction | 72
    acute toxic nephritis | 72
    severe osseous destruction | 72
    superinfection | 72
    below knee amputation rejected | 72
    amputation agreed two weeks later | 72
    surgery performed | 72
    multiorgan dysfunction syndrome | 72
    intensive care efforts | 72
    died | 72
    <|eot_id|>
    