33 years old | 0
unmarried | 0
nullipara | 0
family history of testicular cancer | 0
nonspecific abdominal pain | -1680
explorative laparoscopy | -1680
gelatinous tumor spread detected | -1680
biopsy | -1680
diagnosis of disseminated peritoneal adenomucinosis | -1680
perforated mucinous cystadenoma of the appendix | -1680
advised to undergo peritonectomy and bilateral oophorectomy | -1680
referred for consultation on fertility preservation options | -1680
decided to undergo IVF and embryo cryopreservation | -1680
oocytes retrieved | -1680
embryos fertilized with donor sperm | -1680
embryos cryopreserved | -1680
PMP surgery | 0
extended spread of the disease found | 0
parietal peritoneum resected | 0
omentectomy | 0
appendectomy | 0
splenectomy | 0
bilateral adnexectomy | 0
uterus left intact | 0
postoperatively received heated intraperitoneal infusions of mitomycin C | 0
disease relapsed | 432
elevation of carcinoembrionic antigen | 432
intra abdominal fluid accumulation | 432
multiple peritoneal lesions | 432
explorative laparotomy | 432
cytoreduction and peritonectomy | 432
intraperitoneal infusion of 5-fluorouracil | 432
disease-free for more than 7 years | 8760
desired to become pregnant | 8760
consultation with institutional oncologists | 8760
preparation of the endometrium | 8760
administration of E2 valerate | 8760
vaginal administration of micronized progesterone | 8760
endometrial thickness reached 8 mm | 8760
thawed embryos transferred | 8760
hCG positive | 8760
hCG doubled | 8760
diagnosed with deep vein thrombosis | 1008
started on enoxaparin | 1008
difficult to anatomically identify the uterine cervix on ultrasonography | 1344
urinary bladder appeared to be "smeared" all over the uterus | 1344
left flank pain | 1560
elevation of creatinine | 1560
Betametasone given for fetal lung maturation | 1560
mild bilateral hydronephrosis | 1560
no evidence of urine jets | 1560
urinary bladder covered the anterior part of the uterus | 1560
Doppler USG ruled out renal vein thrombosis | 1560
cystoscopy revealed distorted bladder trigone | 1560
pigtail inserted into the left ureter | 1560
symptoms gradually resolved | 1560
urosepsis | 1680
intravenous antibiotic treatment | 1680
condition improved | 1680
left flank pain | 1792
difficulty in urinating | 1792
blood creatinine sharply risen | 1792
nephrostomy suggested | 1792
decided to deliver the fetus | 1792
oxytocin to induce labor | 1792
vaginal delivery | 1792
healthy male neonate delivered | 1792
transferred to neonatal intensive care unit | 1792
postpartum hemorrhage | 1792
received packed cells | 1792
postpartum course uneventful | 1792
blood creatinine level returned to normal | 1792
put on warfarin | 1792
discharged home | 1792
referred to oncologist, hematologist, and urologist | 1792