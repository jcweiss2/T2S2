66 years old | 0
male | 0
hypertension | 0
hyperlipidemia | 0
hepatitis C virus infection | 0
atrial fibrillation | 0
anticoagulated with apixaban | 0
admitted to the hospital | 0
dizziness | -2
lost consciousness | -2
found down by a family member | -2
Glasgow Coma Score of 15 | 0
no focal neurological deficits | 0
noncontrast CT of the head | 0
right frontal subdural hematoma | 0
right medial orbital wall fracture | 0
no operative intervention recommended | 0
severe headache | 48
head CT repeated | 48
worsening of the subdural hematoma | 48
mass effect | 48
midline shift | 48
no surgical intervention recommended | 48
discharged to acute inpatient rehabilitation | 144
repeat head CT | 216
terrible headache | 216
repeat neurosurgical evaluation | 216
expansion of the hematoma | 216
increased mass effect | 216
midline shift | 216
burr holes for evacuation of the subdural hematoma | 216
placement of subdural drain | 216
headache improved | 222
subdural hematoma decreased in size | 222
drain removed | 222
discharged home | 222
seizure prophylaxis with levetiracetam | 222
strange sensation in the right arm | 338
feeling of inability to control the arm | 338
sent to the emergency room | 338
focal left arm seizure | 338
treated for seizure | 338
started on electroencephalography (EEG) monitoring | 338
admitted | 338
unresponsive | 344
CT head showed no acute hemorrhage | 344
EEG indicated status epilepticus | 344
intubated for airway protection | 344
transferred to the medical intensive care unit | 344
cerebral CTA obtained | 344
negative for any pathology | 344
ventilator-dependent respiratory failure | 344
septic shock secondary to Pseudomonas bacteremia | 344
tracheostomy | 344
gastrostomy | 344
stabilized and discharged to long-term acute care hospital | 413
levetiracetam and oxcarbazepine for seizure control | 413
less responsive | 417
transferred back for neurosurgical evaluation | 417
opened eyes to stimulation | 417
localized with the right upper extremity | 417
minimal movement of left upper and bilateral lower extremities | 417
cough, gag, corneal, and pupillary reflexes were all present | 417
CT and CTA head showed right frontal intraparenchymal hemorrhage | 417
no vascular lesion or anomaly | 417
cerebral catheter angiography performed | 417
prominence of the anterior temporal branch of the right middle cerebral artery | 417
early, rapid, shunting of blood through a cortical vein to the superior sagittal sinus | 417
opacification of a capillary-like serpiginous tangle of vessels | 417
representing an AVM | 417
Spetzler-Martin Grade 1 (Spetzler-Ponce Grade A) | 417
embolization of the AVM performed using N-butyl-cyanoacrylate glue | 425
embolization was successful | 425
no opacification of the early draining vein or AVM nidus | 425
resection of the AVM | 441
right pterional craniotomy performed | 441
AVM separated from surrounding brain parenchyma using microdissection techniques | 441
feeding arteries coagulated using bipolar electrocautery and resected | 441
draining vein coagulated using bipolar electrocautery and resected | 441
intraparenchymal hematoma evacuated | 441
intraoperative Doppler ultrasound indicated no arterial flow in the draining vein | 441
postoperative angiography showed no residual AVM | 441
mental status progressively improved | 449
followed commands and tracked with his eyes | 449
spontaneous antigravity movement of the right upper extremity | 449
no movement of the left upper or bilateral lower extremities | 449
postoperative course complicated by pseudomonas sepsis | 449
treated in consultation with infectious disease | 449
discharged to long-term acute care | 465