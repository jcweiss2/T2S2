44 years old | 0
    male | 0
    Darier6White disease | -8760
    symptom onset during infancy | -43800
    first diagnosed in 1995 | -216576
    mild acne | -43800
    seborrheic distribution | -43800
    summertime exacerbations | -43800
    treated with systemic retinoids | -216576
    multiple complications from 1995 to 2014 | -216576
    sepsis episodes | -216576
    Kaposi varicelliform eruption | -216576
    frequent local infections | -216576
    Staphylococcus aureus infections | -216576
    Morganella morganii infections | -216576
    atypical Mycobacterium cutaneous infection in 2005 | -131040
    infections treated with antibiotics | -216576
    disease peak during 2013 | -17520
    widespread erythema | -17520
    hypertrophic warty keratotic papules | -17520
    plaques | -17520
    cysts | -17520
    nodules | -17520
    giant comedones | -17520
    severe macerations | -17520
    severe fetor | -17520
    leonine-like facies | -17520
    diffuse palmo-plantar keratoderma | -17520
    extreme cachexia | -17520
    tachycardia | -17520
    normal neuropsychiatric evaluation | -17520
    skin biopsy findings | -17520
    keratotic plugs | -17520
    dyskeratosis | -17520
    corps ronds | -17520
    grains | -17520
    suprabasal clefts | -17520
    Periodic acid-Schiff staining negative | -17520
    anemia | -17520
    leukocytosis | -17520
    hypoalbuminemia | -17520
    Staphylococcus aureus skin culture | -17520
    Morganella morganii skin culture | -17520
    Streptococcus group G skin culture | -17520
    S aureus blood culture | -17520
    negative fungal infection tests | -17520
    negative HIV serology | -17520
    negative herpes simplex PCR | -17520
    negative varicella zoster PCR | -17520
    low blood iron | -17520
    low folic acid | -17520
    low transferrin | -17520
    low vitamin D | -17520
    normal immune function tests | -17520
    negative genetic test for 3-base deletion | -17520
    treated with broad-spectrum antibiotics | -17520
    high-dose oral isotretinoin | -17520
    topical keratolytic therapy | -17520
    infections responded well | -17520
    partial response of cutaneous disease | -17520
    discharged | -17520
    presented to ICU 10 months later | -240
    severe sepsis | -240
    severe hypoglycemia | -240
    widespread erythema | -240
    died 2 days after admission | 48

Alright, let's tackle this case report and extract the clinical events with their respective timestamps. 

First, the patient is a 44-year-old male with a unique severe form of Darier2White disease (DWD). The case report mentions that his symptom onset was during infancy, which is around 44 years ago. Since the admission event is at time 0, the symptom onset would be at -44 years, which converts to -44 * 8760 hours/year = -385,440 hours. But wait, the case report says "symptom onset was during infancy" and specifies that mild acne was present since 6 months of age. So, 6 months old is 0.5 years, so 0.5 * 8760 = -4380 hours. Hmm, maybe I need to adjust that.

Wait, the report mentions that the disease was first diagnosed in 1995 when the patient was 27. Since he's 44 now, that means 44 - 27 = 17 years ago. So 17 years * 8760 hours/year = -149,160 hours. But the case report says "data regarding symptoms during infancy were not available, yet according to the patient, mild acne was present in a seborrheic distribution since 6 months of age..." So 6 months is 0.5 years, which is 0.5 * 8760 = -4380 hours. But how does that fit into the timeline?

The first diagnosis in 1995 (17 years ago) would be at -149,160 hours. The symptoms (mild acne, seborrheic distribution, summertime exacerbations) started at 6 months of age, which is 44 years ago minus 6 months? Wait, the patient is 44 now, so 44 years ago is when he was born. 6 months of age would be 43.5 years ago, so 43.5 * 8760 = -381,060 hours. But the admission is at time 0, so all events before admission are negative.

But in the example given earlier, the admission is at 0, and events before have negative times. So the events here: symptom onset during infancy (6 months old) would be -43.5 years converted to hours: -43.5 * 8760 = -381,060 hours. But that seems too far back. The case report says he was first diagnosed in 1995 when he was 27. So 44 - 27 = 17 years ago. So diagnosis in 1995 is -17 * 8760 = -149,160 hours. Then, from 1995 to 2014, he had multiple complications, which would be between -149,160 and - (44-2014) wait, 2014 is 10 years ago (44 now, so 2014 was when he was 34, 44-34=10 years ago). So 10 years ago is -87,600 hours. Wait, maybe I need to adjust the timeline.

Wait, the case report says he was first diagnosed in 1995 at age 27. He is now 44, so 44 - 27 = 17 years since diagnosis. So the diagnosis was 17 years ago, which is -17 * 8760 = -149,160 hours. The complications from 1995 to 2014 (which is a 19-year period from 1995 to 2014) but since he was 27 in 1995 and 44 in the current year, 2014 would be 10 years ago (44 - 34 = 10 years ago). So events from 1995 to 2014 span from -149,160 hours (17 years ago) to -87,600 hours (10 years ago). So the complications during this period would have varying timestamps. But the case report states "from 1995 to 2014 suffered multiple complications including several episodes of sepsis..." So each event in this period would have different timestamps. However, since the exact dates aren't provided, except for the atypical Mycobacterium infection in 2005, which is 2005. If he was 27 in 1995, then in 2005 he was 37, so 44 - 37 = 7 years ago, which is -61,320 hours. 

But the report mentions "an atypical Mycobacterium cutaneous infection in 2005", which is 2005. So 44 now, 2005 was 19 years ago (assuming current year is 2024), so 19 years * 8760 = -166,440 hours. Wait, but the patient's age is 44 now, and the case report was published in 2024? Hmm, the case report's date isn't given, but since the patient is 44 and the last event is death 2 days after admission, which is at +48 hours. So admission is time 0, death at +48.

The key events to extract include:

- Darier-White disease (DWD) diagnosis in 1995 (-149,160 hours)
# 2023-24-project
## This is the project title
### This is a subtitle

This is a paragraph where you can type full text.
You can make *italic* text, **bold** text, or ***combined***.
You can also highlight `code` with backticks.

```python
def hello_world():
  print("Hello World!")
hello_world()
```

```C
#include <stdio.h>
int main(){
  printf("Hello World!");
  return 0;
}
```
[This is a link](https://github.com)

| Header 1 | Header 2 |
|----------|----------|
| Item 1   | Item 2   |
| Item 3   | Item 4   |

- List item 1
Duy
- List item 2
Duy 2
