74 years old | 0
male | 0
admitted to the hospital | 0
unconscious | 0
intubation | 0
hemodynamic stabilization | 0
transferred to cardiac intensive care unit | 0
presumed devastating cardiac event | 0
reactive airway disease | -672
Karo syrup with ephedrine (Forcalide syrup) | -672
ingestion of gasoline | -672
accidental ingestion of gasoline at age 7 | -75936
symptoms of airway disease worsened | -336
doubled daily intake of Karol-Ephedrine syrup | -336
respiratory system improved | -168
returned to usual daily activities | -168
dull epigastric pain | -168
periodic bouts of extreme pain | -168
fever | -168
anorexia | -168
disoriented | -24
febrile | -24
constant extreme abdominal pain | -24
septic shock | 0
abdominal source | 0
rigid and markedly distended abdomen | 0
severe episodes of epigastric pain | 0
massively dilated stomach | 0
decompressed loops of small bowel | 0
nasogastric tube placed | 0
rush of air and 200 ml of blood-stained bilious fluid | 0
exploratory laparotomy | 24
more than 3 liters of transudative ascites evacuated | 24
stomach decompressed | 24
extensive necrosis | 24
multiple microperforations | 24
subtotal gastrectomy | 24
intestinal continuity restored with Roux-en-Y cardiojejunostomy | 24
discharged from the hospital | 168
discontinued use of Karol-Ephedrine syrup | 168
no complications associated with gastrointestinal ischemia | 168
investigated cause of patient's unusual isolated gastric ischemia | 168
sample of Karol-Ephedrine syrup tested | 168
sample of patient's serum tested | 168
ephedrine found in Karol-Ephedrine syrup and serum | 168
hematoxylin and eosin staining of gastrectomy specimen | 168
chronic gastritis | 168
microvascular thrombosis | 168
full thickness necrosis | 168
multiple gastric perforations | 168