65 years old | 0
relapsed ovarian cancer | 0
treated with carboplatin | 0
412 mg dose of carboplatin | 0
dose calculated using Calvert formula | 0
dyspnea | 20
wheezing | 20
hypotension | 20
confusion | 20
blood pressure 90/40 mm Hg | 20
saturation 78% in room air | 20
pulse rate 140 bpm | 20
breath rate 34 breaths/min | 20
infusion stopped | 20
transferred to intensive care unit | 20
intubated | 20
respiratory failure | 20
adrenaline infused | 20
fluids infused | 20
corticosteroids infused | 20
cardiac ultrasound performed | 20
acute coronary syndrome excluded by ECG | 20
acute coronary syndrome excluded by troponin I | 20
pulmonary embolism ruled out by spiral CT scan | 20
Swan-Ganz catheter inserted via right subclavian vein | 20
pulmonary capillary wedge pressure 4 mm Hg | 20
central venous pressure 3 mm Hg | 20
ventilated based on acute respiratory distress syndrome ventilation protocol | 20
blood cultures negative | 20
urine cultures negative | 20
rapid abdomen ultrasound normal | 20
brain CT scan without findings | 20
fever | 168
ventilator-associated pneumonia | 168
bronchoalveolar lavage drawn | 168
treated with antibiotics | 168
became septic | 168
died | unknown
- 65 years old | 0
" relapsed ovarian cancer | 0" (since it's the reason for treatment)
" treated with carboplatin | 0" (as part of the admission)
" 412 mg dose of carboplatin | 0"
" dose calculated using Calvert formula | 0"
blood pressure 90/40 | 20
saturation 78% | 20
pulse 140 | 20
breath rate 34 | 20
transferred to ICU | 20
pulmonary embolism ruled out by CT | 20
Swan-Ganz catheter inserted | 20
ventilated per ARDS protocol | 20
abdomen ultrasound normal | 20
brain CT normal | 20
fever | 164
ventilator-associated pneumonia | 164
bronchoalveolar lavage | 164
treated with antibiotics | 164
became septic | 164 (or later? It says 'thereafter', so maybe after antibiotics, so 164 + some time, but exact time not given, so approximated as 164)
died | unknown (time not specified, so left as unknown)
