70 years old|0
female|0
hypertension|0
hyperlipidaemia|0
diabetes|0
supraventricular tachycardia|0
syncope|-48
weakness|-48
polyuria|-48
elevated blood glucose|-48
negative RT-PCR swab for COVID-19|0
prophylactic anticoagulation|0
transthoracic echocardiogram showing dilated right ventricle|24
computed tomography pulmonary angiogram|48
repeat echocardiogram showing pulmonary embolism and clot in transit|48
therapeutic anticoagulation|48
positive RT-PCR swab for COVID-19|48
percutaneous aspiration thrombectomy with AngioVac|48
death|48
denied fever|0
denied chills|0
denied sore throat|0
denied cough|0
denied chest pain|0
denied dyspnoea|0
initial blood pressure 84/55 mmHg|0
pulse 72 bpm|0
oxygen saturation 88% on room air|0
respiratory rate 16/min|0
temperature 36.6°C|0
no jugular venous distension|0
normal heart sounds|0
normal lung sounds|0
no peripheral edema|0
admitted to telemetry|0
hydration|0
insulin|0
antibiotics|0
droplet precautions|0
contact isolation|0
differential diagnosis: hypovolemia due to diabetic ketoacidosis and sepsis|0
differential diagnosis: acute PE|0
differential diagnosis: myocardial infarction|0
differential diagnosis: arrhythmia|0
differential diagnosis: heart failure|0
suspected underlying COVID-19|0
unremarkable chest X-ray|0
unremarkable head computed tomography|0
electrocardiogram showed sinus rhythm at 80 bpm with S1, Q3, T3 pattern, prolonged QTc, and T-wave inversions across the precordium|0
hyperglycemia (580 mg/dL)|0
elevated anion gap|0
serum creatinine 1.6 mg/dL|0
lactate 7.5 mmol/L|0
D-dimer 2153 ng/mL|0
C-reactive protein 8.6 mg/L|0
pro-BNP 14042 pg/mL|0
INR 1.2|0
negative serial troponin T-tests|0
urine positive for ketones|0
urine positive for white cells|0
blood gas (venous) pH 7.41, pCO2 35.6 mmHg, pO2 30.5 mmHg, HCO3 22 mmol/L, sO2 59.3%|0
white-cell count 14.3 per nL|0
hemoglobin 13.7 g/dL|0
platelet count 210 per nL|0
fibrinogen 182 mg/dL|48
ferritin 61 μg/L|48
procalcitonin NA|48
dyspnea|24
desaturation (93% on 3L oxygen)|24
pulse 80 bpm|24
blood pressure 132/78 mmHg|24
transferred to intensive care unit|48
multidisciplinary institutional PERT evaluation|48
percutaneous aspiration thrombectomy with adjunctive intra-pulmonary and catheter-directed thrombolysis|48
administration of intra-pulmonary and systemic thrombolysis|48
patient arrested|48
