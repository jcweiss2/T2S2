38 years old | 0
woman | 0
admitted to the hospital | 0
fever | -48
nausea | -48
severe sepsis | 0
MSSA bacteraemia | 0
right-sided CRT-D device infection | 0
intravenous antibiotics started | 0
vancomycin | 0
piperacillin-tazobactam | 0
cefazolin monotherapy | 0
transesophageal echocardiogram | 0
no vegetations | 0
device generator extraction | 24
lead extraction | 24
infected pocket debridement | 24
cultures of device generator | 24
cultures of ventricular leads | 24
MSSA growth | 24
suspected endocarditis | 0
normotensive | 0
asymptomatic | 0
AF with complete heart block | 0
junctional escape rhythm | 0
heart rate 40–60 beats per minute | 0
temporary transvenous pacing deferred | 0
transcutaneous pacer pads | 0
dopamine available | 0
blood cultures cleared | 216
no growth | 216
replacement device generator placement | 432
new subxiphoid pocket | 432
biventricular epicardial leads | 432
transthoracic echocardiogram | 432
trivial pericardial effusion | 432
nausea | 504
dizziness | 504
diaphoresis | 504
malaise | 504
blood pressure 79/47 mmHg | 504
paced heart rate 60 beats/min | 504
respiratory rate 20 breaths/min | 504
oxygen saturation 98% | 504
clear breath sounds | 504
elevated jugular venous pressure | 504
distant heart sounds | 504
no rubs | 504
no murmurs | 504
trace pedal pitting edema | 504
pretibial pitting edema | 504
elevated leukocyte count | 504
up-trending leukocyte count | 504
stable hemoglobin | 504
high-sensitivity troponin T flat trend | 504
elevated C-reactive protein | 504
elevated erythrocyte sedimentation rate | 504
normal anti-nuclear antibody | 504
normal C3 complement | 504
normal C4 complement | 504
normal thyroid-stimulating hormone | 504
AF with complete heart block | 504
100% ventricular pacing | 504
enlarged cardiac silhouette | 504
large pericardial effusion | 504
right ventricular collapse | 504
LVEF 30–35% | 504
moderate to large pericardial effusion | 504
diastolic RV collapse | 504
systolic right atrial collapse | 504
lactated ringer's bolus | 504
pericardiocentesis | 504
1L fluid removal | 504
pericardial drain placement | 504
normalized blood pressure | 504
serous fluid analysis | 504
normal nucleated cell count | 504
neutrophilic predominance | 504
pericardial fluid protein 5.6 g/dL | 504
serum protein 5.5 g/dL | 504
no bacterial growth | 504
no fungal growth | 504
colchicine started | 504
chest CT scan | 504
epicardial electrodes in place | 504
pericardial drain output ceased | 672
drain removed | 672
nausea | 672
hypotension | 672
blood pressure 85/59 mmHg | 672
re-accumulation of pericardial effusion | 672
early systolic RA invagination | 672
late diastolic RV collapse | 672
repeat pericardiocentesis | 672
1.5L fluid removal | 672
pericardial drain placement | 672
prednisone added | 672
ibuprofen added | 672
transthoracic echocardiogram | 672
increased pericardial effusion size | 672
no tamponade signs | 672
transthoracic pleuro-pericardial window | 744
small-bore chest tube placement | 744
drainage decline | 744
transthoracic echocardiogram | 912
no significant pericardial effusion | 912
discharged home | 912
chest tube in place | 912
colchicine continued | 912
ibuprofen continued | 912
prednisone taper | 912
intravenous cefazolin continued | 912
stable at 1-month follow-up | 1344
asymptomatic | 1344
minimal chest tube drainage | 1344
repeat TTE at 2 months | 1440
no effusion | 1440
chest tube removed | 1440
repeat TTE at 4 months | 2928
no effusion | 2928
feeling well | 2928
