29 years old | 0
male | 0
admitted to the hospital | 0
breathlessness | -336
cough with white sputum | -168
loss of weight and appetite | -420
shooting pain in the right side of chest | -168
blood pressure of 110/70 | 0
respiratory rate of 28/min | 0
oxygen saturation (SpO2) of 90% on room air | 0
cardiomegaly | 0
pleural effusion with fissural extension | 0
underlying collapse on the right side with fibrotic bands in right perihilar region | 0
Total leucocyte count (TLC) count was 10,730 cells | 0
neutrophilic predominance | 0
pleural tap of 300 ml fluid | 0
exudative effusion | 0
intercostal drain (ICD) insertion | 0
diagnosis of lower respiratory tract infection | 0
treated with intravenous antibiotics | 0
nebulizations | 0
other supportive measures | 0
pleural fluid analysis | 0
sugars 75 mg/dl | 0
proteins <2 g/dl | 0
adenosine deaminase (ADA) 4.8 u/l | 0
pleural fluid cytology | 0
white blood cells of 950 cells | 0
lymphocytic (95%) | 0
reactive mesothelial cells | 0
left atrial wall thickening | 0
infiltration or thrombus | 0
pulmonary vein obstruction | 0
good left ventricle function | 0
homogeneous poorly enhancing soft tissue in subcarinal region | 0
indenting left atrium | 0
partial narrowing of right inferior pulmonary vein ostium | 0
extending along the interatrial groove | 0
encasing mass | 0
partial narrowing of the right main pulmonary artery | 0
azygous arch | 0
cervical mediastinoscopy and biopsy of 4R lymph node station | 0
frozen section was remained inconclusive | 0
discharged | 120
underwent VATS and incisional biopsy | 168
hard mass encasing heart and hilar structures | 168
infiltrating left atrium | 168
biopsy for histopathological examination and immunohistochemistry | 168
extubated | 168
received noninvasive ventilation and oxygen (O2) support | 168
developed tachypnea | 192
shifted back to surgical intensive care unit | 192
procalcitonin levels were raised | 192
D-dimer levels were within normal limits | 192
arterial blood gas showed partial pressure 54.5 | 192
SpO2 of 90% on bilevel positive airway pressure with O2 support of 10 L | 192
intubated | 192
connected to ventilator support | 192
ET culture and sensitivity | 192
Gram stain | 192
fungal stain | 192
acid-fast bacilli stain | 192
ET culture sensitivity | 192
Gram-negative coverage | 192
X-ray postintubation showed left lower lobe pneumonia | 192
basal crept bilaterally | 192
blood culture was negative | 192
endotracheal secretion culture grown pseudo hyphae | 192
hyaline septate with acute branching hyphae | 192
started on voriconazole 200mg BID therapy | 192
HPE report revealed several epithelioid granulomas | 192
numerous multinucleated giant cells | 192
areas of necrotising inflammation | 192
few scattered acute branching fungal hyphae | 192
diagnosis of acute respiratory distress syndrome with invasive aspergillosis | 192
treated accordingly with low tidal volume strategy | 192
condition worsened | 216
developed septic shock | 216
refractory hypoxemia | 216
serum creatinine increased to 3.1 mg/dl | 216
developing acute kidney injury | 216
started on renal replacement therapy | 216
hyperkalemia | 216
acidosis | 216
family refused to take any further treatment | 216
left against medical advice | 216
expired | 216
cardiac arrest | 216