51 years old | 0
male | 0
admitted to the hospital | 0
right chest and back pain | -720
no family and other medical history | 0
biopsy | -720
needle aspiration | -720
diagnose the right lower pulmonary pseudotumor | -720
wedge resection of the right lower lobe | -720
CT scan | 0
mass in the lower lobe of the right lung | 0
bone destruction of the 7, 8, and 9 thoracic vertebrae | 0
multiple enlarged lymph nodes | 0
bilateral pleural hypertrophy | 0
fibre cord signs | 0
informed consent | 0
general anesthesia | 7
thoracic vertebral lesions removed | 7
right lung lesions | 7
needle aspiration | 7
pathological examination | 7
acute and chronic purulent inflammations | 7
inflammatory granulation and granuloma | 7
tuberculosis could not be excluded | 7
sputum culture | 7
negative | 7
postoperative pathological consultations | 7
neutrophils, lymphocytes, monocytes, scattered eosinophils, multinucleated giant-cell infiltration, and fibrinous exudation | 7
fibrinous exudation | 7
organization in the alveolar cavity | 7
neutrophils, lymphocytes, monocytes, scattered multinucleated giant-cell infiltration, and significant focal necrosis | 7
necrosis | 7
neutrophil aggregation and abscesses | 7
special infectious disease | 7
non-caseating necrosis | 7
neutrophil aggregation | 7
abscesses | 7
Department of Hematology | 7
bone biopsy | 7
increased plasma cells | 7
myeloma could not be excluded | 7
high fever | 24
antibiotics and antipyretic treatment | 24
improved | 24
left upper arm was painful | 672
CT imaging | 672
destruction in the 8th to 10th ribs | 672
malignant tumors suspected | 672
pleural effusion | 672
solitary nodule | 672
malignant tumors suspected | 672
striped high-density shadows | 672
inflammatory lesions | 672
multiple enlarged lymph nodes | 672
malignant bone tumors | 672
left humeral tumor lesion removal | 720
osteoma-like hyperplasia | 720
hemorrhaging | 720
inflammatory granulation tissues and granulomas | 720
pus samples | 720
drug sensitivity tests | 720
no bacterial growth | 720
postoperative CT scan | 744
peripheral lung cancer | 744
inflammatory pseudotumor | 744
prednisone acetate tablets | 744
oral | 744
30 mg/day | 744
6 weeks | 744
reduced | 744
percutaneous puncture biopsy | 816
argon-helium knife ablation | 816
CT scans | 816
puncture needle | 816
tissue | 816
knives | 816
treatment | 816
local edema | 816
bleeding | 816
chronic inflammation | 816
fibrous tissues | 816
inflammatory granulation tissue | 816
compound cyclophosphamide tablets | 1008
50 mg/day | 1008
2 weeks | 1008
discontinued | 1008
bone marrow suppression | 1008
hemoglobin | 1008
91 g/L | 1008
71 g/L | 1008
shortness of breath | 1008
improved | 1008
discharged | 1008
admitted to hospital for the 2nd time | 1344
chest CT scan | 1344
left upper lobe nodules | 1344
enlarged | 1344
patched high-density shadows | 1344
observed | 1344
lung inflammatory pseudotumor | 1344
benign | 1344
malignant tendency | 1344
severe pain | 1344
radiation therapy | 1368
20 Gy/10 F | 1368
re-examination of chest CT scans | 1404
left upper lobe nodule | 1404
right lung lamella | 1404
smaller | 1404
shadow | 1404
lighter | 1404
admitted to hospital for the 3rd time | 2160
severe anemia | 2160
red-blood cell transfusion | 2160
nutritional support | 2160
symptomatic treatment | 2160
hematological consultation | 2160
recombinant human granulocyte colony stimulating factor | 2160
rhGCSF | 2160
promote bone marrow erythroid hematopoiesis | 2160
anti-infection | 2160
phlegm treatments | 2160
pulmonary infection | 2160
anemia | 2160
improved | 2160
discharged | 2304
admitted to hospital for the 4th time | 2880
aggravated left humerus pain | 2880
MRI | 2880
chronic osteomyelitis | 2880
peripheral inflammatory pseudotumor | 2880
infection | 2880
routine antibiotic treatment | 2880
poor effect | 2880
debridement | 2912
osteomyelitis | 2912
soft tissue infection | 2912
pathological diagnosis | 2912
inflammatory granulation tissues | 2912
granuloma | 2912
purulent necrosis | 2912
supportive treatments | 2912
lung infection | 2912
urinary tract infection | 2912
sputum culture | 2912
urine culture | 2912
antimicrobial susceptibility tests | 2912
antibiotic therapy | 2912
condition | 2912
improved | 2912
discharged | 2976
admitted to hospital for the 5th time | 3504
breathing difficulties | 3504
unconsciousness | 3504
Orthopedics Department | 3504
severe pneumonia | 3504
septic shock | 3504
multiple organ dysfunction syndromes | 3504
metabolic acidosis | 3504
type II respiratory failure | 3504
osteomyelitis | 3504
soft tissue infection | 3504
urinary system infection | 3504
hypoalbuminemia | 3504
incomplete paralysis | 3504
postoperative right pulmonary pseudotumor | 3504
increasing chest tightness | 3504
intensive care unit | 3504
anti-infection | 3504
anti-inflammatory | 3504
expectorant | 3504
electrolyte imbalance | 3504
condition | 3504
not improved | 3504
active treatment | 3504
ceased | 3504
died | 3504
septic shock | 3504
cause of death | 3504
no autopsy | 3504