69 years old | 0
male | 0
admitted to the hospital | 0
chronic weakness | -8760
recurrent admissions | -8760
untreated and undiagnosed pancytopenia | -8760
splenomegaly | -8760
neutropenia | -8760
fungal pneumonia | -720
aspergilloma | -720
Pneumocystis jirovecii pneumonia | -720
right thyroidectomy | -8760
thyroid cancer | -8760
posterior right coronary artery stenting | -8760
chronic stable angina pectoris | -8760
paroxysmal atrial fibrillation | -8760
exacerbation of fungal pneumonia | 0
afebrile | 0
body temperature 36.5°C | 0
blood pressure 99/66 mm Hg | 0
heart rate 77 beats per minute | 0
respiratory rate 20 per minute | 0
poor nutritional status | 0
weight 48.7 kg | 0
height 169 cm | 0
body mass index 17.05 kg/m2 | 0
cachectic | 0
exhausted | 0
pancytopenia | 0
neutropenia | 0
hyponatremia | 0
increased prothrombin time | 0
increased partial thromboplastin time | 0
elevated C-reactive protein | 0
elevated erythrocyte sedimentation rate | 0
no evidence of cytomegalovirus infection | 0
no other causes of atypical pneumonia | 0
negative blood cultures | 0
negative sputum cultures | 0
urine culture positive for Gram-positive cocci | 0
multiple nodular consolidations in the left upper lung | 0
multiple nodular consolidations in the right upper lobe | 0
left pleural effusion | 0
pericardial effusion | 0
no enlarged lymph nodes | 0
enlarged spleen | 0
aspirin | 0
nicorandil | 0
trimetazidine | 0
bisoprolol | 0
levothyroxine | 0
total parenteral nutrition | 0
antibiotic therapy | 0
trimethoprim/sulfamethoxazole | 0
meropenem | 0
amphotericin B | 0
cefepime | 0
consultations from hematology | 0
consultations from rheumatology | 0
consultations from infection | 0
differential diagnosis | 0
splenomegaly | 0
normochromic normocytic anemia | 0
reticulocyte percentage 0.65% | 0
anemia of chronic disease | 0
elevated ferritin | 0
low transferrin | 0
normal serum iron level | 0
no deficiency of B12 and folate | 0
bone marrow biopsy | 0
average cellularity 60% | 0
no signs of bone marrow failure | 0
positive anti-nuclear antibodies | 0
rheumatoid factor | 0
weakly-positive anti-DNA | 0
anti-cardiolipin immunoglobulin M antibodies | 0
low serum C3 | 0
normal C4 | 0
oral ulcer | 0
no other autoimmune features | 0
elevated cystatin C | 0
cystatin C-based estimated glomerular filtration rate 42.6 mL/min/1.73 m2 | 0
normal creatinine level | 0
indeterminate renal function | 0
equivocal levels of anti-DNA antibodies | 24
splenectomy | 240
partial splenic embolization | 384
infusion of 1.5 L of fluid | 264
transfusion of filtered red blood cells | 264
norepinephrine | 264
sepsis | 264
body temperature 37.0°C | 264
blood pressure 86/52 mm Hg | 264
pulse rate 84 | 264
partial splenic embolization | 384
iodixanol | 384
ultrasound guidance | 384
right common femoral artery | 384
celiac angiography | 384
splenic angiography | 384
gelfoam | 384
increase in blood counts | 408
white blood cell count 820/μL | 408
hemoglobin 10.0 g/dL | 408
platelet count 45×103/μL | 408
temperature 38.5°C | 432
decrease in blood pressure to 84/56 mm Hg | 432
pulse rate increase to 148 per minute | 432
septic shock | 432
norepinephrine and fluids | 432
CT scans of the chest and abdomen | 432
no pulmonary embolism | 432
no bowel perforation | 432
mechanical ventilation | 456
cardiac arrest | 480
cardiopulmonary resuscitation | 480
death | 480