56 years old | 0
male | 0
ST-elevation myocardial infarction | 0
transported to the catheterization lab | 0
primary percutaneous intervention | 0
left anterior descending artery occlusion | 0
thrombus aspiration | 0
stent implementation | 0
no-reflow phenomenon | 0
hemodynamic instability | 0
ventricular fibrillation | 0
pulseless electrical activity | 0
CPR commenced | 0
LUCAS3™ device use | 0
decision to use ECMO | 0
2 rounds of CPR | 0
no return of spontaneous circulation | 0
cannulation | 0
hemodynamic improvement | 0
CPR discontinued | 0
PCI finished | 0
LAD flow restored | 0
three-vessel disease | 0
transported to ICU | 0
ECMO support | 0
waking up | 24
mechanical ventilation weaned | 24
no significant neurological consequences | 24
deterioration | 24
lactate 15.3 mmol/l | 24
high doses of vasopressors | 24
high doses of inotropes | 24
norepinephrine 0.36 mcg/kg/min | 24
terlipressin 0.67 mcg/kg/min | 24
adrenaline 0.21 mcg/kg/min | 24
cannula positions checked | 24
X-ray | 24
ultrasound | 24
ECMO machine operating appropriately | 24
hemoglobin fall from 14.5 g/dl to 8.3 g/dl | 24
suspected bleeding in right proximal leg or pelvis | 24
repeated attempts to achieve distal perfusion | 24
local hematoma | 24
massive blood transfusion protocol | 24
packed red blood cells 15 units | 24
fresh frozen plasma 3 units | 24
cryoprecipitate 10 units | 24
platelets 20 units | 24
lactate dropped to 6 mmol/l | 24
hemoglobin raised to 11.2 g/dl | 24
short-term improvement | 24
abdominal compartment syndrome | 48
inflated abdomen | 48
intraabdominal hypertension 16 cmH2O | 48
declining urine output | 48
creatinine 2.6 mg/dl | 48
increased vasopressor doses | 48
lactate raised to 14 mmol/l | 48
hemoglobin not improved beyond 11 g/dl | 48
PRBC rapid infusions 2 | 48
transported for abdominal CT | 72
significant hemoperitoneum | 72
grade IV liver lacerations | 72
consultation with general surgeons | 72
transported to operating room | 72
general anesthesia | 72
left lobectomy | 72
extubated | 96
condition improved | 96
vasopressors reduced | 96
lactate levels normalized | 96
PRBC transfusions 3 | 96
hemoglobin maintained at 10-11 g/dl | 96
second echocardiogram | 168
ejection fraction improved to 30-35% | 168
considered for ECMO weaning | 168
arrhythmias | 192
non-sustained ventricular tachycardia | 192
ventricular fibrillation | 192
defibrillations | 192
repeat echocardiography | 216
ejection fraction reduced to 16% | 216
arrhythmias stabilized | 216
decision to transfer for LVAD implantation | 216
transferred to another hospital | 216
ECMO support | 216
spontaneous breathing with nasal prongs | 216
hemodynamic stability | 216
no vasopressors | 216
awake | 216
alert | 216
no gross neurological sequelae | 216
catastrophic multiorgan failure | 264
sepsis | 264
death | 264
