65 years old|0
    female|0
    rheumatic valve disease|0
    surgical mitral valve repair|0
    percutaneous exchange of the mitral valve|0
    dyspnea on the slightest effort|0
    paroxysmal nocturnal dyspnea|0
    orthopnea|0
    dry cough|0
    daily episodes of fever between 38 and 38.5 °C|0
    treated for dengue fever|-960
    episode of paroxysmal atrial flutter|0
    decreased level of consciousness (Glasgow coma scale of 13)|0
    anisocoric pupils|0
    referred to the intensive care unit (ICU)|0
    drowsy|0
    pale|0
    hydrated|0
    acyanotic|0
    anicteric|0
    afebrile (37.3 °C)|0
    arterial blood pressure 122/73 mm Hg|0
    heart rate 96 beats per minute|0
    respiratory rate 14 breaths per minute|0
    heart auscultation normal|0
    murmurs absent|0
    respiratory auscultation normal|0
    abdomen examination normal|0
    mild edema in the lower limbs|0
    hemoglobin 8.5 g/dL|0
    hematocrit 25%|0
    white blood cells 16,200/mm³|0
    platelets 192,000/mm³|0
    no left shift|0
    mild anisocytosis|0
    microcytosis|0
    urea 67 mg/dL|0
    creatinine 2.39 mg/dL|0
    sodium 132 mmol/L|0
    potassium 3.6 mmol/L|0
    C reactive protein 11.2 mg/dL|0
    APACHE II score 22 (death risk 45%)|0
    SAPS III score 64 (death risk 44%)|0
    precarious dentition|0
    blood culture samples collected|0
    empirical treatment with ceftriaxone|0
    gentamicin initiated|0
    transesophageal echocardiogram revealed vegetation|0
    decreased level of consciousness|240
    sensitive conduction aphasia|240
    mild right central paralysis|240
    ischemic stroke suspected|240
    brain tomography demonstrated hypodense left insular lobe|240
    mechanical thrombectomy indicated|240
    arteriogram did not show occlusion of proximal vessels|240
    failed partial filling of the parietal branch of the left middle cerebral artery|240
    worsened level of consciousness|240
    hemodynamic instability|240
    need for hemodialysis|240
    orotracheal intubation performed|240
    vasoactive drugs initiated|240
    repeated brain tomography|240
    brain edema in the posterior circulation region|240
    hypodensity in the left thalamus|240
    septic shock refractory to therapeutic measures|240
    died|240
    transesophageal echocardiogram showed left atrial dilation|0
    moderate double mitral lesion|0
    mild to moderate tricuspid insufficiency|0
    moderate pulmonary hypertension|0
    vegetation confirmed|0
    Haemophilus parainfluenzae in blood cultures|0
    sensitive to B-lactamic compounds|0
    systemic embolism suspected|0
    central nervous system involvement|240
    middle cerebral artery affected|240
    pulmonary embolism risk|240
    abscess formation risk|240
    severe valve dysfunction risk|240
    chordae rupture risk|240
    early identification of etiological agent|0
    empirical antibiotic use|0
    high sensitivity to penicillin|0
    high sensitivity to cephalosporins|0
    early administration of antimicrobial|0
    difficulty isolating Haemophilus parainfluenzae|0
    
    65 years old|0
    female|0
    rheumatic valve disease|0
    surgical mitral valve repair|0
    percutaneous exchange of the mitral valve|0
    dyspnea on the slightest effort|0
    paroxysmal nocturnal dyspnea|0
    orthopnea|0
    dry cough|0
    daily episodes of fever between 38 and 38.5 °C|0
    treated for dengue fever|-960
    episode of paroxysmal atrial flutter|0
    decreased level of consciousness (Glasgow coma scale of 13)|0
    anisocoric pupils|0
    referred to the intensive care unit (ICU)|0
    drowsy|0
    pale|0
    hydrated|0
    acyanotic|0
    anicteric|0
    afebrile (37.3 °C)|0
    arterial blood pressure 122/73 mm Hg|0
    heart rate 96 beats per minute|0
    respiratory rate 14 breaths per minute|0
    heart auscultation normal|0
    murmurs absent|0
    respiratory auscultation normal|0
    abdomen examination normal|0
    mild edema in the lower limbs|0
    hemoglobin 8.5 g/dL|0
    hematocrit 25%|0
    white blood cells 16,200/mm³|0
    platelets 192,000/mm³|0
    no left shift|0
    mild anisocytosis|0
    microcytosis|0
    urea 67 mg/dL|0
    creatinine 2.39 mg/dL|0
    sodium 132 mmol/L|0
    potassium 3.6 mmol/L|0
    C reactive protein 11.2 mg/dL|0
    APACHE II score 22 (death risk 45%)|0
    SAPS III score 64 (death risk 44%)|0
    precarious dentition|0
    blood culture samples collected|0
    empirical treatment with ceftriaxone|0
    gentamicin initiated|0
    transesophageal echocardiogram revealed vegetation|0
    decreased level of consciousness|240
    sensitive conduction aphasia|240
    mild right central paralysis|240
    ischemic stroke suspected|240
    brain tomography demonstrated hypodense left insular lobe|240
    mechanical thrombectomy indicated|240
    arteriogram did not show occlusion of proximal vessels|240
    failed partial filling of the parietal branch of the left middle cerebral artery|240
    worsened level of consciousness|240
    hemodynamic instability|240
    need for hemodialysis|240
    orotracheal intubation performed|240
    vasoactive drugs initiated|240
    repeated brain tomography|240
    brain edema in the posterior circulation region|240
    hypodensity in the left thalamus|240
    septic shock refractory to therapeutic measures|240
    died|240
    transesophageal echocardiogram showed left atrial dilation|0
    moderate double mitral lesion|0
    mild to moderate tricuspid insufficiency|0
    moderate pulmonary hypertension|0
    vegetation confirmed|0
    Haemophilus parainfluenzae in blood cultures|0
    sensitive to B-lactamic compounds|0
    systemic embolism suspected|240
    central nervous system involvement|240
    middle cerebral artery affected|240
    pulmonary embolism risk|240
    abscess formation risk|240
    severe valve dysfunction risk|240
    chordae rupture risk|240
    early identification of etiological agent|0
    empirical antibiotic use|0
    high sensitivity to penicillin|0
    high sensitivity to cephalosporins|0
    early administration of antimicrobial|0
    difficulty isolating Haemophilus parainfluenzae|0