23 years old | 0
multipara | 0
admitted to the Intensive Care Unit | 0
spontaneous vaginal delivery | -48
live full-term male baby | -48
hemodynamic instability | 0
febrile | 48
severe abdominal pain | 48
lower abdominal quadrant pain | 48
elevated D-dimer | 48
elevated C-reactive protein | 48
received cefazoline | 48
received low molecular weight heparin | 48
hypotensive | 48
aggressive fluid resuscitation | 48
contrast-enhanced computerized tomography | 48
thrombus in one of the right pelvic veins | 48
dilated right ureter | 48
dilated right renal pelvis | 48
elevated procalcitonin | 48
elevated urea | 48
elevated creatinine | 48
metronidazole added to therapy | 48
transferred to ICU | 48
vasopressors not needed | 48
antibiotic therapy changed | 48
ceftriaxone used | 48
dosage of LMWH increased | 48
episodes of tachypnea | 72
peaks of body temperature elevation | 72
falls in peripheral oxygen saturation | 72
hypoxemia | 72
hypocapnia | 72
pulmonary congestion | 72
bilateral parenchymal infiltrates | 72
pleural effusion | 72
intensive respiratory physiotherapy | 72
noninvasive ventilation | 72
conventional mechanical ventilation not needed | 72
microbiological cultures negative | 72
cervical smear revealed Streptococcus pyogenes group A | 72
transferred to High Dependency Unit | 72
antibiotic therapy with metronidazole discontinued | 168
LMWH discontinued | 168
dismissed for home care | 336
referred to hematologist | 336