63 years old | 0
male | 0
admitted to the hospital | 0
signet ring cell carcinoma | -672
neoadjuvant chemotherapy | -672
gastrectomy | -672
Roux-en-Y reconstruction | -672
infrarenal AAA | -504
diameter of AAA 4.1 cm | -504
follow-up | -504
admitted to the hospital | 0
urosepsis | 0
pyelonephritis | 0
anaemia | 0
Hb 85 g/L | 0
WBC 33.3 × 10^9/L | 0
CRP 87 mg/L | 0
PCT 3.3 ng/mL | 0
CTA scan | 0
AAA enlargement | 0
thrombosed intramural haematoma | 0
subfebrile fever | 240
constipation | 240
severe fatigue | 240
anaemia | 240
Hb 78 g/L | 240
Hct 23% | 240
CRP 123 g/L | 240
PCT 6.5 ng/mL | 240
negative faecal occult blood test | 240
absent GI tract bleeding symptoms | 240
ruptured AAA | 240
pseudoaneurysm | 240
urgent operation | 240
total laparotomy | 240
enlarged pulsating inflammatory conglomerate | 240
PAEF | 240
duodenal compression | 240
necrotic pars ascendens | 240
infrarenal cross-clamping technique | 240
resection of infrarenal AAA | 240
replacement with Dacron graft | 240
resection of pars horizontalis and pars ascendens | 240
postoperative recovery | 240
readmitted to the hospital | 2880
recurrent fainting episodes | 2880
pain in the abdomen | 2880
haematemesis | 2880
severe idiopathic hypoglycaemia | 2880
RBC transfusions | 2880
CT scans | 2880
gastroscopies | 2880
coloscopies | 2880
capsule-endoscopy | 2880
jejunal ulcer | 2880
PET scan | 2880
metabolically active regions | 2880
total laparotomy | 2880
SAEF | 2880
defect in the jejunum | 2880
infrarenal aortic cross-clamping | 2880
removal of Dacron graft | 2880
replacement with xenograft | 2880
intravenous antibiotic therapy | 2880
per os acetylsalicylic acid | 2880
follow-up CTA | 4320
patent aortic graft | 4320
no signs of inflammation or fistulisation | 4320