29 years old | 0
    African American | 0
    male | 0
    SCD (Hb SS) | 0
    exchange transfusions every 4-6 wk | 0
    hemosiderosis | 0
    cirrhosis | 0
    vaso-occlusive pain crisis in lower extremities | 0
    uncontrolled epistaxis | 0
    deferasirox | 0
    folic acid | 0
    oxycodone | 0
    denied tobacco | 0
    denied alcohol | 0
    denied drug use | 0
    jaundiced | 0
    alert | 0
    fully oriented | 0
    soft abdomen | 0
    no tenderness | 0
    no organomegaly | 0
    normal bowel sounds | 0
    new-onset confusion | 24
    hepatic encephalopathy | 24
    conjugated hyperbilirubinemia | 0
    total serum bilirubin 57 mg/dL | 0
    direct serum bilirubin 30 mg/dL | 0
    alkaline phosphatase 306 U/L | 0
    aspartate transaminase 227 U/L | 0
    alanine transaminase 54 U/L | 0
    white blood cell count 38.6 k/µL | 0
    hemoglobin 6.3 g/dL | 0
    platelet count 39 k/µL | 0
    negative Coomb's testing | 0
    fibrinogen 412 mg/dL | 0
    INR 2.3 | 0
    MELD-sodium score 40 | 0
    acute liver injury | 0
    negative viral hepatitis testing | 0
    negative autoimmune hepatitis testing | 0
    negative genetic testing | 0
    ferritin 1399 ng/mL | 0
    arterial ammonia 72 µmol/L | 0
    acute kidney injury | 0
    serum creatinine 3.48 mg/dL | 0
    cirrhosis | 0
    patent hepatic vasculature | 0
    normal hepatic flow | 0
    no biliary ductal dilatation | 0
    acute-on-chronic liver failure | 0
    multi-system organ failure | 0
    acute sickle cell intrahepatic cholestasis | 0
    new-onset acute liver injury | 0
    encephalopathy | 0
    coagulopathy | 0
    admitted to medical intensive liver unit | 0
    intubation | 0
    mechanical ventilation | 0
    acute hypoxic respiratory failure | 0
    acute chest syndrome | 0
    vancomycin | 0
    meropenem | 0
    exchange transfusion initiated | 0
    HbS decrease from 56.3 to 8.2 g/dL | 0
    no improvement in hepatic synthetic function | 0
    listed for urgent liver transplantation | 0
    pre-operative evaluation | 0
    multidisciplinary team involvement | 0
    underwent liver transplantation | 216
    standard piggyback technique | 216
    duct-to-duct biliary anastomosis | 216
    enlarged explanted liver | 216
    focally micronodular capsule | 216
    congested parenchyma | 216
    normal hepatic vasculature | 216
    normal bile ducts | 216
    sinusoidal dilatation | 216
    sickled RBC clusters | 216
    pigmented histiocytes | 216
    cholestasis | 216
    sinusoidal fibrosis | 216
    portal-portal bridging fibrosis | 216
    cirrhosis | 216
    hepatocellular siderosis | 216
    Kupffer cell siderosis | 216
    exchange transfusion resumed | 216
    immunosuppression induction therapy | 216
    antithymocyte globulin | 216
    mycophenolate mofetil | 216
    tacrolimus | 216
    steroid taper | 216
    HCV RNA >100000000 IU/mL | 216
    HCV genotype 1A | 216
    glecaprevir/pibrentasvir started | 552
    discharged | 552
    sustained virologic response | 3240
    preserved liver synthetic function | 8760
    monthly exchange transfusions | 8760
    target HbS <20% | 8760

    