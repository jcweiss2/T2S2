23 years old | 0
male | 0
deceased-donor renal transplant | -12000
end-stage renal disease | -12000
membranoproliferative glomerulonephritis | -12000
tacrolimus | -12000
prednisone | -12000
fever | -336
fatigue | -336
intermittent fever | -336
intermittent fatigue | -336
admitted to the hospital | 0
blood pressure 112/67 mmHg | 0
heart rate 103 beats per minute | 0
pulse oximetry 98% | 0
temperature 37.1°C | 0
body mass index 22.6 kg/m² | 0
S3 | 0
holosystolic murmur | 0
scattered crackles | 0
mild peripheral edema | 0
coronavirus 2019 PCR testing negative | 0
borderline sinus tachycardia | 0
pulmonary edema | 0
leukocytosis | 0
thrombocytosis | 0
mild acute kidney injury | 0
elevated cardiac troponin | 0
elevated NT-prohormone-brain natriuretic peptide | 0
elevated D-dimer | 0
hospitalized | 0
meropenem | 0
linezolid | 0
levofloxacin | 0
fluconazole | 0
low-dose nitroglycerin | 0
furosemide infusions | 0
vegetation on the anterior mitral valve leaflet | 0
perforation | 0
ruptured chordae tendinae | 0
torrential mitral regurgitation | 0
Coandă effect | 0
vegetation on the aortic valve | 0
torrential aortic regurgitation | 0
infectious diseases team consulted | 24
serology testing | 24
Bartonella henselae antibody IgM positive | 24
Bartonella henselae antibody IgG positive | 24
Coxiella burnetii phase I IgM antibodies positive | 24
Coxiella burnetii phase I IgG antibodies positive | 24
Coxiella burnetii phase II IgM antibodies positive | 24
Coxiella burnetii phase II IgG antibodies positive | 24
doxycycline | 24
gentamicin | 24
transesophageal echocardiography | 72
bicuspid aortic valve | 72
dual valve replacement | 168
aspirin | 168
warfarin | 168
international normalized ratio 2.5 | 168
outpatient clinics | 240
hydroxychloroquine therapy | 720
clinically well | 2160
no prosthetic valve endocarditis | 2160
no valve dysfunction | 2160