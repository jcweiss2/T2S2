34 years old | 0 | 0 
male | 0 | 0 
primary refractory acute myeloblastic leukemia | -8760 | -8760 
allogeneic bone marrow transplant | -648 | -648 
delayed engraftment | -648 | 0 
prolonged severe neutropenia | -648 | 0 
vancomycin-resistant Enterococcus | -648 | 0 
Streptococcus viridans | -648 | 0 
Streptococcus mitis | -648 | 0 
bacteremia | -648 | 0 
tedizolid | -648 | 0 
cefepime | -648 | 0 
Flagyl | -648 | 0 
daptomycin | -648 | 0 
filgrastim | 0 | 0 
acyclovir | 0 | 0 
Bactrim | 0 | 0 
caspofungin | 0 | 0 
acute abdominal pain | 0 | 0 
fever | 0 | 0 
tachycardia | 0 | 0 
hypotension | 0 | 0 
tachypnea | 0 | 0 
distended abdomen | 0 | 0 
localized peritonitis | 0 | 0 
white cell count 0.2 x 10^9 /L | 0 | 0 
absolute neutrophil count (ANC) of zero | 0 | 0 
anemic | 0 | 0 
hemoglobin of 7 g/L | 0 | 0 
thrombocytopenic | 0 | 0 
platelet count of 10 x 10^9 /L | 0 | 0 
lactic acid of 3.1 mmol/L | 0 | 0 
CT scan | 0 | 0 
segmental ischemia of the small bowel | 0 | 0 
exploratory laparotomy | 0 | 24 
ischemic bowel segment | 0 | 24 
small bowel resection | 0 | 24 
primary anastomosis | 0 | 24 
norepinephrine | 0 | 24 
vasopressin | 0 | 24 
transesophageal echo | 0 | 24 
intensive care unit | 24 | 48 
pressors weaned | 24 | 48 
extubated | 48 | 48 
transferred to the floor | 48 | 48 
diet advanced | 72 | 72 
passed flatus | 72 | 72 
new fevers | 96 | 96 
increased abdominal pain | 96 | 96 
lactic acidosis | 96 | 96 
respiratory decompensation | 96 | 96 
neutropenic | 96 | 96 
white cell count of 0.1 x 10^9 /L | 96 | 96 
ANC 0 | 96 | 96 
lactic acid 3.7 mmol/L | 96 | 96 
amphotericin B | 96 | 120 
repeat CT scan | 96 | 120 
necrotic small bowel | 96 | 120 
expedited pathology report | 96 | 120 
invasive fungal forms | 96 | 120 
omental and small intestinal resection specimens | 96 | 120 
hematologic dissemination of mucormycosis | 96 | 120 
septic emboli | 96 | 120 
comfort measures | 120 | 120 
died | 120 | 120 
mucormycosis | -648 | 120 
angioinvasion | -648 | 120 
vessel thrombosis | -648 | 120 
tissue necrosis | -648 | 120 
disseminated | -648 | 120 
rhinocerebral | -648 | 120 
pulmonary | -648 | 120 
cutaneous | -648 | 120 
gastrointestinal systems | -648 | 120 
colon | -648 | 120 
diagnosis | -648 | 120 
culture | -648 | 120 
histopathology | -648 | 120 
serum fungal tests | -648 | 120 
1,3-beta-D-glucan | -648 | 120 
Aspergillus galactomannan | -648 | 120 
PCR | -648 | 120 
amphotericin B lipid complex | -648 | 120 
posaconazole | -648 | 120 
surgical debulking | -648 | 120 
typhlitis | -648 | 120 
hemodynamic instability | -648 | 120 
left lower quadrant pain | 0 | 0 
expeditious surgical resection | 0 | 24 
antifungal coverage | 0 | 120 
amphotericin | 96 | 120 
repeat exploratory laparotomy | 120 | 120 
bowel resection | 120 | 120 
prognosis | 120 | 120