37 years old | 0
female | 0
admitted to the hospital | 0
altered mental state | 0
cortisol-secreting ACC | -540
adrenalectomy | -540
recurrent lesion | -270
radical nephrectomy | -270
adjuvant radiotherapy | -270
hypercortisolemia | -180
chemotherapy with Avastin + FOLFOX | -30
mental change | 0
septic shock | 0
respiratory failure | 0
fluid resuscitation | 0
vasopressor support | 0
invasive ventilation | 0
white blood cell count = 140/mm3 | 0
hemoglobin level = 7.2 g/dL | 0
platelet count = 8,000/mm3 | 0
total bilirubin level = 1.6 mg/dl | 0
serum aspartate aminotransferase/alanine aminotransferase = 102/102 IU/L | 0
blood urea nitrogen/serum creatinine = 24.1/1.12 mg/dL | 0
lactic acid level = 8.13 mmol/L | 0
c-reactive protein level = 21.86 mg/dl | 0
procalcitonin level = 42.46 ng/ml | 0
lobar consolidation in the right lower lung zone (RLLZ) | 0
neutropenic septic shock | 0
pneumonia | 0
catheter-related infection | 0
antibiotics (meropenem, vancomycin) | 0
central catheter removal | 0
vasopressor taper | 24
mechanical ventilation discontinuation | 96
neutrophil count recovery | 72
MRSA identified | 48
septic shock relapse | 120
respiratory failure relapse | 120
re-intubation | 120
multifocal ground-glass opacities | 120
elevated serum galactomannan titer | 120
Aspergillus fumigatus growth | 120
intravenous voriconazole | 120
P. jirovecii observed | 120
pneumocystis pneumonia diagnosis | 120
trimethoprim/sulfamethoxazole | 120
MRSA bacteremia persistence | 120
vancomycin to linezolid switch | 168
Candida albicans growth | 168
candidemia resolution | 168
combined bacterial pneumonia | 168
mitotane therapy | 168
cortisol level decrease | 168
hemoptysis | 240
pneumonia-associated cavitary lesion | 240
ventilator readings deterioration | 240
oxygen requirements increase | 240
peritoneal seeding | 720
lymph node metastases | 720
do-not-resuscitate order | 720
discharge | 720
death | 744