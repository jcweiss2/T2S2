27 years old | 0
    man | 0
    admitted to the hospital | 0
    pancytopenia | 0
    neutrophils: 0.8×109/L | 0
    hemoglobin: 9.4 gr/dl | 0
    platelets: 4×109/L | 0
    muco-cutaneous hemorrhages | 0
    severe aplastic anemia | 0
    empirical broad spectrum antibiotherapy | 120
    piperacillin–tazobactam | 120
    amikacin | 120
    febrile neutropenia | 120
    fever | 120
    fever resolved | 120
    neutropenia worsened | 0.3×109/L | 168
    oral prednisone | 288
    admitted to the intensive care unit | 456
    septic shock | 456
    prednisone stopped | 456
    piperacillin-tazobactam restarted | 480
    levofloxacin | 480
    blood cultures positive | Streptococcus mitis | 480
    blood cultures positive | Klebsiella pneumoniae | 480
    recovered | 576
    admitted to hematology unit | 576
    central venous catheter inserted | 600
    fever reappeared | 696
    piperacillin–tazobactam replaced | meropenem | 696
    levofloxacin replaced | meropenem | 696
    antifungal treatment initiated | caspofungin | 696
    fever persisted | 696
    poor clinical condition | 696
    diarrhea | 696
    abdominal pain | 696
    dry cough | 696
    left thoracic pain | 696
    peripheral blood cultures positive | septate hyphae | 744
    central venous blood cultures positive | septate hyphae | 744
    caspofungin replaced | liposomal amphotericin B | 744
    caspofungin replaced | voriconazole | 744
    stool examination | S. clavata | 528
    CT scan | left pulmonary nodular lesion | 744
    diffuse bowel thickening | 744
    multiple nodular lesions | spleen | 744
    multiple nodular lesions | kidneys | 744
    multiple nodular lesions | liver | 744
    normal liver function tests | 744
    CVC removed | 744
    left blurred vision | 744
    cerebral CT scan normal | 744
    cerebral magnetic resonance imaging normal | 744
    retinal hemorrhage | 744
    echocardiogram excluded fungal endocarditis | 744
    severe neutropenia | <0.1×109/L | 744
    S. clavata identified | blood culture | 792
    clinical condition improved | 792
    daily blood cultures positive | S. clavata | 792
    weekly stool examinations negative | 792
    daily blood cultures negative | 792
    fever persisted | 1008
    no documented infection | 1008
    negative galactomannan antigenemia | 1008
    voriconazole blood levels | 2.4 µg/mL | 1008
    antifungal susceptibility testing | echinocandins | high MICs | 1008
    fluconazole | high MIC | 1008
    amphotericin B | low MIC | 1008
    5-fluorocytosine | low MIC | 1008
    voriconazole | low MIC | 1008
    posaconazole | low MIC | 1008
    allogeneic bone marrow transplantation | 1008
    conditioning regimen | cyclophosphamide | 840
    conditioning regimen | fludarabine | 840
    conditioning regimen | alemtuzumab | 864
    cyclosporine started | 1008
    granulocyte transfusions | days 39, 40, 41, 48, 49 | 936, 960, 984, 1152, 1176
    neutrophil counts | 0.5–1×109/L | post-transfusion
    neutrophil counts | <0.1×109/L | without transfusion
    fever resolved | 1008
    good clinical condition | 1008
    neutrophil count | 0.5×109/L | 1632
    voriconazole replaced by posaconazole | 2016
    nausea and vomiting | 2016
    liposomal amphotericin B discontinued | 2016
    abdominal ultrasound | small splenic residual lesions | 2016
    left hospital | 2112
    posaconazole secondary prophylaxis | 2112
    fever resolved | 2112
    vision normalized | 2112
    no recurrence of infection | 4-month follow-up
    no complications of transplantation | 4-month follow-up