39 years old | 0
female | 0
type 2 diabetes | -672
deep vein thrombosis | -672
gastritis | -672
schizophrenia | -672
self-harm | -672
admitted to the medical admissions unit | 0
right sub-mammary abscess | -168
spreading cellulitis of the breast | -168
septic | 0
pyrexia of 39.2 | 0
blood pressure of 127/65 | 0
tachycardia of 110 | 0
widespread cellulitis involving the nipple and sub-mammary area | 0
cellulitis spreading to the axilla | 0
white cell count of 23.8 | 0
neutrophils 19.9 | 0
CRP of 428 | 0
simple cellulitis diagnosed | 0
commenced on parenteral antibiotics | 0
fluid resuscitation | 0
intravenous benzyl penicillin | 0
flucloxacillin | 0
condition worsened | 72
sought surgical opinion | 72
evidence of synergistic gangrene | 72
cellulitis spread | 72
areas of growing necrotic ulceration | 72
resuscitation commenced | 72
antibiotic therapy adjusted | 72
imipenem | 72
clindamycin | 72
taken to theatre | 75
partial mastectomy performed | 75
wound left open and packed | 75
postoperatively stable on intensive care | 75
returned to theatre for further debridement | 96
radical debridement performed | 96
further debridement performed | 96
wound monitored closely | 120
vacuum dressing applied | 120
signs of sepsis improved | 120
returned to the ward | 120
nutritional supplements | 120
adequate hydration | 120
secondary closure performed | 312
preoperative cultures taken | 75
mixture of gram positive and negative bacteria | 75
Bacteroides spp | 75
sensitive to metronidazole | 75
sensitive to clindamycin | 75
sensitive to imipenem | 75
histology confirmed widespread microscopic changes | 75
abscess formation consistent with gangrene | 75
no evidence of malignancy | 75
blood markers of infection improved | 120
no signs of secondary organ failure | 120
discharged | 528
intravenous antibiotics administered | 75
changed to oral antibiotics | 240
co amoxiclav | 240
metronidazole | 240
follow-up arranged | 528
possibility of reconstruction considered | 528