28 years old | 0
male | 0
admitted to the hospital | 0
burn injuries | -72
intubated | -72
airway protection | -72
minimal ventilatory support | -72
oxygen saturation 100% | 0
arterial partial pressure of oxygen 326 mm Hg | 0
crystalloid fluid resuscitation | 0
Parkland formula | 0
hypoxemia | 72
increased inspired oxygen fraction | 72
high positive end-expiratory pressure | 72
sedated | 72
neuromuscular blockade | 72
Pao2/Fio2 50 mm Hg | 72
pulmonary bilateral infiltrates | 72
ARDS | 72
VV-ECMO | 96
reinfusion cannula placement | 96
drainage cannula placement | 96
ECMO flows 4.7 to 5.0 L/min | 96
Spo2 >90% | 96
oxygenation status worsened | 120
Pao2/Fio2 43 mm Hg | 120
elevated cardiac output | 120
ECMO flow/native CO ratio 0.45 to 0.50 | 120
reconfigured veno-VV-ECMO circuit | 144
increased flows to 6 to 6.5 L/min | 144
hypoxemia not corrected | 144
lactate dehydrogenase elevated | 144
postoxygenator Pao2 100 to 200 mm Hg | 144
second ECMO circuit inserted in parallel | 168
combined flow 6 L/min | 168
ECMO postoxygenator Pao2 >350 mm Hg | 168
patient's Spo2 >90% | 168
lactate dehydrogenase decreased | 168
respiratory status improved | 192
Pao2/Fio2 430 mm Hg | 192
heavy diuresis | 192
pulmonary hygiene | 192
ventilator settings weaned to Fio2 40% | 192
weaned down to one system | 216
weaning process | 216
decreased flows on additional system | 216
patient tolerated single system configuration | 216
weaned off remaining circuit | 240
decannulated completely from ECMO | 240
sepsis | 240
pneumonia | 240
bacteremia | 240
fungemia | 240
gastrointestinal bleeding | 240
multiple debridements | 240
skin grafts | 240
discharged on room air | 720
total hospital stay 3 months | 720