66 years old | 0
male | 0
admitted to the hospital | 0
asthenia | -24
adynamia | -24
mild dyspnoea | -24
dry cough | -24
chills | -24
fever | -24
diaphoresis | -24
altered consciousness state | -24
disorientation | -24
episodes of agitation | -24
great respiratory difficulty | -24
desaturation | -24
hypertensive nephropathy | -8760
polycystic kidney disease | -8760
renal transplantation | -720
immunosuppressive treatment | -720
tacrolimus | -720
prednisolone | -720
azathioprine | -720
chest x-ray | 0
consolidation in the middle third of the left pulmonary field | 0
respiratory failure | 24
invasive mechanical ventilation support | 24
septic shock | 24
multiple organ failure syndrome | 24
neurological compromise | 24
stupor | 24
empirical antibiotic treatment | 24
piperacillin/tazobactam | 24
vancomycin | 24
clarithromycin | 24
fluconazole | 24
oseltamivir | 24
urinary antigen testing for Histoplasma | 48
urinary antigen testing for Cryptococcus | 48
bronchoalveolar lavage galactomannan test | 48
liposomal amphotericin B | 96
ganciclovir | 48
viral load for cytomegalovirus | 48
blood cultures | 48
oral tracheal secretion cultures | 48
brain tomography | 72
intra-axial lesion | 72
ring enhancement | 72
vasogenic oedema | 72
cerebritis | 72
open biopsy | 96
subcortical mass | 96
fresh examination | 96
microbiological studies | 96
histopathological studies | 96
septate dematiaceous hyphae | 96
amphotericin B | 96
voriconazole | 96
neurosurgical intervention | 120
ventilation support discontinued | 120
alertness restored | 120
Sabouraud agar | 120
growth of flat, cottony, grey-white colonies | 120
greenish black colonies | 120
dark brown colour | 120
microbiological typing | 144
phaeohyphomycosis | 144
disseminated Alternaria spp. | 144
MRI scan | 120
collection on the surgical bed | 120
oedema in the right subinsular region | 120
terbinafine treatment | 120
computed tomography scans | 240
no significant changes in brain lesions | 240
no progression of mycosis | 240
no other organs compromised | 240
death | 2880