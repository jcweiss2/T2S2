27 years old | 0
male | 0
ulcerative colitis | -672
primary sclerosing cholangitis | -672
total abdominal colectomy with end-ileostomy | -672
abdominal pain | -168
high ileostomy output | -168
9-kg weight loss | -168
admitted to the Emergency Department | 0
tachycardia | 0
afebrile | 0
blood pressure of 103/74 mm Hg | 0
dilated loops of bowel to the level of the colostomy | 0
white blood cell count of 5.4 K/uL | 0
alanine aminotransferase of 446 unit/L | 0
aspartate aminotransferase of 268 unit/L | 0
alkaline phosphatase of 1034 unit/L | 0
point of care lactate of 3.32 mmol/L | 0
admitted to the ward of colorectal surgery services | 0
nil-per-os status | 0
resuscitated with 1900 mL of intravenous fluids | 0
nasogastric tube was placed | 0
metoprolol tartrate 25 mg twice daily | 0
hydromorphone 0.2 mg every 4 h | 0
ondansetron 4 mg every 6 h | 0
acetaminophen 1000 mg every 8 h | 0
pantoprazole 40 mg | 0
tachycardia | 24
fever | 72
tachypnea | 72
leukopenia | 72
mild agitation | 72
worsening abdominal pain | 72
upgraded to the ICU | 72
IVF resuscitation | 72
broad spectrum antibiotics | 72
piperacillin-tazobactam 3.375 g every 6 h | 72
metoprolol tartrate 12.5 mg | 72
thyroid function testing | 72
thyroid-stimulating hormone levels below detectable limits | 72
elevated levels of triiodothyronine | 72
elevated levels of tetraiodothyronine | 72
normal parathyroid hormone level | 72
diagnosis of hyperthyroidism | 72
diagnosis of thyroid storm | 72
esmolol infusion | 72
propylthiouracil 150 mg every 6 h | 72
cholestyramine 4 mg twice daily | 72
intravenous hydrocortisone 50 mg every 8 h | 72
continuous IVF hydration | 72
acetaminophen 1000 mg as needed | 72
elevated thyroid-stimulating immunoglobulins level | 96
ileostomy output decreased | 96
fevers resolved | 168
discharged home | 408
propranolol 30 mg twice daily | 408
propylthiouracil 200 mg twice daily | 408
prednisone 10 mg | 408