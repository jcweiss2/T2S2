76 years old | 0
male | 0
admitted to the hospital | 0
left knee pain | -96
febrile | 0
Glasgow coma scale of 14/15 | 0
heart rate was 125 bpm | 0
polypneic at 25c/min | 0
swelling measuring 15 cm on the inner side of his left thigh | 0
skin necrosis | 0
inflammatory signs | 0
swelling measuring 5 cm in the left inguinal region | 0
leukocytosis of 30,000E/ml | 0
C-reactive protein of 400 mg/l | 0
computed tomography (CT) angiography | 0
diagnosis of septic shock related to necrotizing fasciitis | 0
necrotizing fasciitis of the left thigh | 0
abdominal wall | 0
operation under general anesthesia | 0
hypotensive | 0
tachycardia at 150 bpm | 0
incision in the left inner thigh | 1
pus removal | 1
dissection into quadriceps muscle plains | 1
drainage of 200 milliliters of pus | 1
necrotic debris excised | 1
incision in the left inguinal region | 2
dissection into muscle plans | 2
drainage of 100 milliliters of pus | 2
abdominal midline incision | 3
tumor in the sigmoid | 3
perforated in the retroperitoneum | 3
colostomy on the left flank | 3
biopsy of the tumor | 3
pathological examination | 4
Lieberkuhnian adenocarcinoma | 4
bacteriological examination | 4
E. coli multi-drug-sensitive | 4
negative anerobic culture | 4
septic shock | 0
deceased | 24
colon cancer | -96 
unresectable tumor | 3 
subcutaneous emphysema | 0 
intraoperative view | 3 
retroperitoneal abscess | -96 
femoral ring | -96 
weight loss | -96 
transit disorders | -96 
abdominal pain | -96 
unexplained soft tissue infections | -96 
urgent CT scans | 0 
aggressive surgical debridement | 1 
intensive support | 1 
intravenous antibiotics | 1 
systemic toxicity | 1 
operative debridement | 1 
necrotic material removal | 1 
defect | 4 
antimicrobial | 1 
surgical debridement | 1 
treatment of NF | 1 
NF diagnosis | 0 
NF treatment | 1 
NF management | 1 
NF clinical presentation | -96 
NF suspicion | -96 
NF diagnosis delay | -96 
NF mortality | 24 
NF incidence | -96 
NF etiology | -96 
NF pathogenesis | -96 
NF clinical features | -96 
NF imaging | 0 
NF surgery | 1 
NF sepsis | 0 
NF septic shock | 0 
NF intensive care | 1 
NF antimicrobial therapy | 1 
NF supportive measures | 1 
NF prognosis | 24 
NF outcome | 24 
NF follow-up | 24 
NF recurrence | 24 
NF complication | 24 
NF comorbidity | -96 
NF risk factor | -96 
NF prevention | -96 
NF education | -96 
NF awareness | -96 
NF research | -96 
NF publication | -96 
NF guideline | -96 
NF protocol | -96 
NF algorithm | -96 
NF decision-making | -96 
NF patient care | 1 
NF patient outcome | 24 
NF patient education | -96 
NF patient awareness | -96 
NF patient empowerment | -96 
NF patient support | -96 
NF family support | -96 
NF healthcare provider | 1 
NF healthcare system | 1 
NF quality of care | 1 
NF quality of life | 24 
NF cost-effectiveness | -96 
NF cost-benefit | -96 
NF resource utilization | 1 
NF resource allocation | -96 
NF policy | -96 
NF legislation | -96 
NF advocacy | -96 
NF ethics | -96 
NF law | -96 
NF malpractice | -96 
NF negligence | -96 
NF liability | -96 
NF standard of care | 1 
NF best practice | 1 
NF evidence-based practice | 1 
NF clinical practice guideline | -96 
NF patient safety | 1 
NF medical error | -96 
NF near miss | -96 
NF adverse event | 24 
NF sentinel event | 24 
NF root cause analysis | -96 
NF quality improvement | -96 
NF patient-centered care | 1 
NF family-centered care | -96 
NF culturally competent care | -96 
NF patient engagement | -96 
NF shared decision-making | -96 
NF informed consent | 0 
NF advance care planning | -96 
NF end-of-life care | 24 
NF palliative care | 24 
NF hospice care | 24 
NF bereavement care | 24 
NF spiritual care | -96 
NF chaplaincy care | -96 
NF social work | -96 
NF case management | -96 
NF care coordination | 1 
NF transition of care | 24 
NF readmission | 24 
NF hospitalization | 0 
NF length of stay | 24 
NF intensive care unit | 1 
NF mechanical ventilation | 1 
NF vasopressor | 1 
NF antibiotic | 1 
NF fluid resuscitation | 1 
NF blood transfusion | -96 
NF surgery complication | 24 
NF surgical site infection | -96 
NF wound care | 1 
NF dressing | 1 
NF wound debridement | 1 
NF negative pressure wound therapy | -96 
NF skin graft | -96 
NF flap reconstruction | -96 
NF amputation | -96 
NF disability | 24 
NF rehabilitation | -96 
NF physical therapy | -96 
NF occupational therapy | -96 
NF speech therapy | -96 
NF cognitive therapy | -96 
NF mental health | -96 
NF anxiety | -96 
NF depression | -96 
NF post-traumatic stress disorder | -96 
NF substance abuse | -96 
NF addiction | -96 
NF withdrawal | -96 
NF delirium | -96 
NF dementia | -96 
NF cognitive impairment | -96 
NF neurological deficit | -96 
NF neuropathy | -96 
NF myopathy | -96 
NF radiculopathy | -96 
NF pain management | 1 
NF pain assessment | 1 
NF pain treatment | 1 
NF opioid | 1 
NF non-opioid | 1 
NF adjuvant therapy | 1 
NF alternative therapy | -96 
NF complementary therapy | -96 
NF integrative therapy | -96 
NF nutrition | 1 
NF hydration | 1 
NF electrolyte management | 1 
NF fluid management | 1 
NF medication management | 1 
NF pharmacotherapy | 1 
NF medication adherence | -96 
NF medication non-adherence | -96 
NF medication error | -96 
NF adverse drug reaction | -96 
NF allergic reaction | -96 
NF anaphylaxis | -96 
NF medication side effect | -96 
NF laboratory test | 0 
NF imaging study | 0 
NF diagnostic test | 0 
NF monitoring | 1 
NF vital sign | 0 
NF hemodynamic monitoring | 1 
NF cardiac monitoring | 1 
NF respiratory monitoring | 1 
NF oxygen saturation | 1 
NF capnography | -96 
NF electroencephalogram | -96 
NF electromyogram | -96 
NF nerve conduction study | -96 
NF pulmonary function test | -96 
NF sleep study | -96 
NF polysomnogram | -96 
NF actigraphy | -96 
NF quality metric | -96 
NF performance measure | -96 
NF benchmarking | -96 
NF quality improvement initiative | -96 
NF patient satisfaction | -96 
NF patient experience | -96 
NF family satisfaction | -96 
NF family experience | -96 
NF staff satisfaction | -96 
NF staff experience | -96 
NF healthcare provider satisfaction | -96 
NF healthcare provider experience | -96 
NF leadership | -96 
NF management | -96 
NF governance | -96 
NF policy development | -96 
NF policy implementation | -96 
NF policy evaluation | -96 
NF accreditation | -96 
NF certification | -96 
NF licensure | -96 
NF credentialing | -96 
NF privileging | -96 
NF peer review | -96 
NF quality assurance | -96 
NF quality control | -96 
NF risk management | -96 
NF patient safety program | -96 
NF patient safety initiative | -96 
NF patient safety goal | -96 
NF patient safety objective | -96 
NF patient safety target | -96 
NF patient safety metric | -96 
NF patient safety measure | -96 
NF patient safety benchmark | -96 
NF patient safety best practice | -96 
NF patient safety guideline | -96 
NF patient safety protocol | -96 
NF patient safety algorithm | -96 
NF patient safety decision-making | -96 
NF patient safety education | -96 
NF patient safety training | -96 
NF patient safety awareness | -96 
NF patient safety empowerment | -96 
NF patient safety support | -96 
NF family safety | -96 
NF family education | -96 
NF family training | -96 
NF family awareness | -96 
NF family empowerment | -96 
NF family support | -96 
NF healthcare provider safety | -96 
NF healthcare provider education | -96 
NF healthcare provider training | -96 
NF healthcare provider awareness | -96 
NF healthcare provider empowerment | -96 
NF healthcare provider support | -96 
NF staff safety | -96 
NF staff education | -96 
NF staff training | -96 
NF staff awareness | -96 
NF staff empowerment | -96 
NF staff support | -96 
NF leadership safety | -96 
NF leadership education | -96 
NF leadership training | -96 
NF leadership awareness | -96 
NF leadership empowerment | -96 
NF leadership support | -96 
NF management safety | -96 
NF management education | -96 
NF management training | -96 
NF management awareness | -96 
NF management empowerment | -96 
NF management support | -96 
NF governance safety | -96 
NF governance education | -96 
NF governance training | -96 
NF governance awareness | -96 
NF governance empowerment | -96 
NF governance support | -96 
NF policy safety | -96 
NF policy education | -96 
NF policy training | -96 
NF policy awareness | -96 
NF policy empowerment | -96 
NF policy support | -96 
NF procedure safety | -96 
NF procedure education | -96 
NF procedure training | -96 
NF procedure awareness | -96 
NF procedure empowerment | -96 
NF procedure support | -96 
NF protocol safety | -96 
NF protocol education | -96 
NF protocol training | -96 
NF protocol awareness | -96 
NF protocol empowerment | -96 
NF protocol support | -96 
NF guideline safety | -96 
NF guideline education | -96 
NF guideline training | -96 
NF guideline awareness | -96 
NF guideline empowerment | -96 
NF guideline support | -96 
NF algorithm safety | -96 
NF algorithm education | -96 
NF algorithm training | -96 
NF algorithm awareness | -96 
NF algorithm empowerment | -96 
NF algorithm support | -96 
NF decision-making safety | -96 
NF decision-making education | -96 
NF decision-making training | -96 
NF decision-making awareness | -96 
NF decision-making empowerment | -96 
NF decision-making support | -96 
NF communication safety | -96 
NF communication education | -96 
NF communication training | -96 
NF communication awareness | -96 
NF communication empowerment | -96 
NF communication support | -96 
NF teamwork safety | -96 
NF teamwork education | -96 
NF teamwork training | -96 
NF teamwork awareness | -96 
NF teamwork empowerment | -96 
NF teamwork support | -96 
NF handoff safety | -96 
NF handoff education | -96 
NF handoff training | -96 
NF handoff awareness | -96 
NF handoff empowerment | -96 
NF handoff support | -96 
NF transition safety | -96 
NF transition education | -96 
NF transition training | -96 
NF transition awareness | -96 
NF transition empowerment | -96 
NF transition support | -96 
NF discharge safety | -96 
NF discharge education | -96 
NF discharge training | -96 
NF discharge awareness | -96 
NF discharge empowerment | -96 
NF discharge support | -96 
NF readmission safety | -96 
NF readmission education | -96 
NF readmission training | -96 
NF readmission awareness | -96 
NF readmission empowerment | -96 
NF readmission support | -96 
NF hospital-acquired condition | -96 
NF hospital-acquired infection | -96 
NF central line-associated bloodstream infection | -96 
NF catheter-associated urinary tract infection | -96 
NF ventilator-associated pneumonia | -96 
NF surgical site infection | -96 
NF pressure ulcer | -96 
NF fall | -96 
NF medication error | -96 
NF adverse drug reaction | -96 
NF allergic reaction | -96 
NF anaphylaxis | -96 
NF sentinel event | -96 
NF near miss | -96 
NF adverse event | -96 
NF root cause analysis | -96 
NF quality improvement initiative | -96 
NF patient safety initiative | -96 
NF patient safety goal | -96 
NF patient safety objective | -96 
NF patient safety target | -96 
NF patient safety metric | -96 
NF patient safety measure | -96 
NF patient safety benchmark | -96 
NF patient safety best practice | -96 
NF patient safety guideline | -96 
NF patient safety protocol | -96 
NF patient safety algorithm | -96 
NF patient safety decision-making | -96 
NF patient safety education | -96 
NF patient safety training | -96 
NF patient safety awareness | -96 
NF patient safety empowerment | -96 
NF patient safety support | -96 
NF family safety | -96 
NF family education | -96 
NF family training | -96 
NF family awareness | -96 
NF family empowerment | -96 
NF family support | -96 
NF healthcare provider safety | -96 
NF healthcare provider education | -96 
NF healthcare provider training | -96 
NF healthcare provider awareness | -96 
NF healthcare provider empowerment | -96 
NF healthcare provider support | -96 
NF staff safety | -96 
NF staff education | -96 
NF staff training | -96 
NF staff awareness | -96 
NF staff empowerment | -96 
NF staff support | -96 
NF leadership safety | -96 
NF leadership education | -96 
NF leadership training | -96 
NF leadership awareness | -96 
NF leadership empowerment | -96 
NF leadership support | -96 
NF management safety | -96 
NF management education | -96 
NF management training | -96 
NF management awareness | -96 
NF management empowerment | -96 
NF management support | -96 
NF governance safety | -96 
NF governance education | -96 
NF governance training | -96 
NF governance awareness | -96 
NF governance empowerment | -96 
NF governance support | -96 
NF policy safety | -96 
NF policy education | -96 
NF policy training | -96 
NF policy awareness | -96 
NF policy empowerment | -96 
NF policy support | -96 
NF procedure safety | -96 
NF procedure education | -96 
NF procedure training | -96 
NF procedure awareness | -96 
NF procedure empowerment | -96 
NF procedure support | -96 
NF protocol safety | -96 
NF protocol education | -96 
NF protocol training | -96 
NF protocol awareness | -96 
NF protocol empowerment | -96 
NF protocol support | -96 
NF guideline safety | -96 
NF guideline education | -96 
NF guideline training | -96 
NF guideline awareness | -96 
NF guideline empowerment | -96 
NF guideline support | -96 
NF algorithm safety | -96 
NF algorithm education | -96 
NF algorithm training | -96 
NF algorithm awareness | -96 
NF algorithm empowerment | -96 
NF algorithm support | -96 
NF decision-making safety | -96 
NF decision-making education | -96 
NF decision-making training | -96 
NF decision-making awareness | -96 
NF decision-making empowerment | -96 
NF decision-making support | -96 
NF communication safety | -96 
NF communication education | -96 
NF communication training | -96 
NF communication awareness | -96 
NF communication empowerment | -96 
NF communication support | -96 
NF teamwork safety | -96 
NF teamwork education | -96 
NF teamwork training | -96 
NF teamwork awareness | -96 
NF teamwork empowerment | -96 
NF teamwork support | -96 
NF handoff safety | -96 
NF handoff education | -96 
NF handoff training | -96 
NF handoff awareness | -96 
NF handoff empowerment | -96 
NF handoff support | -96 
NF transition safety | -96 
NF transition education | -96 
NF transition training | -96 
NF transition awareness | -96 
NF transition empowerment | -96 
NF transition support | -96 
NF discharge safety | -96 
NF discharge education | -96 
NF discharge training | -96 
NF discharge awareness | -96 
NF discharge empowerment | -96 
NF discharge support | -96 
NF readmission safety | -96 
NF readmission education | -96 
NF readmission training | -96 
NF readmission awareness | -96 
NF readmission empowerment | -96 
NF readmission support | -96 
NF hospital-acquired condition | -96 
NF hospital-acquired infection | -96 
NF central line-associated bloodstream infection | -96 
NF catheter-associated urinary tract infection | -96 
NF ventilator-associated pneumonia | -96 
NF surgical site infection | -96 
NF pressure ulcer | -96 
NF fall | -96 
NF medication error | -96 
NF adverse drug reaction | -96 
NF allergic reaction | -96 
NF anaphylaxis | -96 
NF sentinel event | -96 
NF near miss | -96 
NF adverse event | -96 
NF root cause analysis | -96 
NF quality improvement initiative | -96 
NF patient safety initiative | -96 
NF patient safety goal | -96 
NF patient safety objective | -96 
NF patient safety target | -96 
NF patient safety metric | -96 
NF patient safety measure | -96 
NF patient safety benchmark | -96 
NF patient safety best practice | -96 
NF patient safety guideline | -96 
NF patient safety protocol | -96 
NF patient safety algorithm | -96 
NF patient safety decision-making | -96 
NF patient safety education | -96 
NF patient safety training | -96 
NF patient safety awareness | -96 
NF patient safety empowerment | -96 
NF patient safety support | -96 
NF family safety | -96 
NF family education | -96 
NF family training | -96 
NF family awareness | -96 
NF family empowerment | -96 
NF family support | -96 
NF healthcare provider safety | -96 
NF healthcare provider education | -96 
NF healthcare provider training | -96 
NF healthcare provider awareness | -96 
NF healthcare provider empowerment | -96 
NF healthcare provider support | -96 
NF staff safety | -96 
NF staff education | -96 
NF staff training | -96 
NF staff awareness | -96 
NF staff empowerment | -96 
NF staff support | -96 
NF leadership safety | -96 
NF leadership education | -96 
NF leadership training | -96 
NF leadership awareness | -96 
NF leadership empowerment | -96 
NF leadership support | -96 
NF management safety | -96 
NF management education | -96 
NF management training | -96 
NF management awareness | -96 
NF management empowerment | -96 
NF management support | -96 
NF governance safety | -96 
NF governance education | -96 
NF governance training | -96 
NF governance awareness | -96 
NF governance empowerment | -96 
NF governance support | -96 
NF policy safety | -96 
NF policy education | -96 
NF policy training | -96 
NF policy awareness | -96 
NF policy empowerment | -96 
NF policy support | -96 
NF procedure safety | -96 
NF procedure education | -96 
NF procedure training | -96 
NF procedure awareness | -96 
NF procedure empowerment | -96 
NF procedure support | -96 
NF protocol safety | -96 
NF protocol education | -96 
NF protocol training | -96 
NF protocol awareness | -96 
NF protocol empowerment | -96 
NF protocol support | -96 
NF guideline safety | -96 
NF guideline education | -96 
NF guideline training | -96 
NF guideline awareness | -96 
NF guideline empowerment | -96 
NF guideline support | -96 
NF algorithm safety | -96 
NF algorithm education | -96 
NF algorithm training | -96 
NF algorithm awareness | -96 
NF algorithm empowerment | -96 
NF algorithm support | -96 
NF decision-making safety | -96 
NF decision-making education | -96 
NF decision-making training | -96 
NF decision-making awareness | -96 
NF decision-making empowerment | -96 
NF decision-making support | -96 
NF communication safety | -96 
NF communication education | -96 
NF communication training | -96 
NF communication awareness | -96 
NF communication empowerment | -96 
NF communication support | -96 
NF teamwork safety | -96 
NF teamwork education | -96 
NF teamwork training | -96 
NF teamwork awareness | -96 
NF teamwork empowerment | -96 
NF teamwork support | -96 
NF handoff safety | -96 
NF handoff education | -96 
NF handoff training | -96 
NF handoff awareness | -96 
NF handoff empowerment | -96 
NF handoff support | -96 
NF transition safety | -96 
NF transition education | -96 
NF transition training | -96 
NF transition awareness | -96 
NF transition empowerment | -96 
NF transition support | -96 
NF discharge safety | -96 
NF discharge education | -96 
NF discharge training | -96 
NF discharge awareness | -96 
NF discharge empowerment | -96 
NF discharge support | -96 
NF readmission safety | -96 
NF readmission education | -96 
NF readmission training | -96 
NF readmission awareness | -96 
NF readmission empowerment | -96 
NF readmission support | -96 
NF hospital-acquired condition | -96 
NF hospital-acquired infection | -96 
NF central line-associated bloodstream infection | -96 
NF catheter-associated urinary tract infection | -96 
NF ventilator-associated pneumonia | -96 
NF surgical site infection | -96 
NF pressure ulcer | -96 
NF fall | -96 
NF medication error | -96 
NF adverse drug reaction | -96 
NF allergic reaction | -96 
NF anaphylaxis | -96 
NF sentinel event | -96 
NF near miss | -96 
NF adverse event | -96 
NF root cause analysis | -96 
NF quality improvement initiative | -96 
NF patient safety initiative | -96 
NF patient safety goal | -96 
NF patient safety objective | -96 
NF patient safety target | -96 
NF patient safety metric | -96 
NF patient safety measure | -96 
NF patient safety benchmark | -96 
NF patient safety best practice | -96 
NF patient safety guideline | -96 
NF patient safety protocol | -96 
NF patient safety algorithm | -96 
NF patient safety decision-making | -96 
NF patient safety education | -96 
NF patient safety training | -96 
NF patient safety awareness | -96 
NF patient safety empowerment | -96 
NF patient safety support | -96 
NF family safety | -96 
NF family education | -96 
NF family training | -96 
NF family awareness | -96 
NF family empowerment | -96 
NF family support | -96 
NF healthcare provider safety | -96 
NF healthcare provider education | -96 
NF healthcare provider training | -96 
NF healthcare provider awareness | -96 
NF healthcare provider empowerment | -96 
NF healthcare provider support | -96 
NF staff safety | -96 
NF staff education | -96 
NF staff training | -96 
NF staff awareness | -96 
NF staff empowerment | -96 
NF staff support | -96 
NF leadership safety | -96 
NF leadership education | -96 
NF leadership training | -96 
NF leadership awareness | -96 
NF leadership empowerment | -96 
NF leadership support | -96 
NF management safety | -96 
NF management education | -96 
NF management training | -96 
NF management awareness | -96 
NF management empowerment | -96 
NF management support | -96 
NF governance safety | -96 
NF governance education | -96 
NF governance training | -96 
NF governance awareness | -96 
NF governance empowerment | -96 
NF governance support | -96 
NF policy safety | -96 
NF policy education | -96 
NF policy training | -96 
NF policy awareness | -96 
NF policy empowerment | -96 
NF policy support | -96 
NF procedure safety | -96 
NF procedure education | -96 
NF procedure training | -96 
NF procedure awareness | -96 
NF procedure empowerment | -96 
NF procedure support | -96 
NF protocol safety | -96 
NF protocol education | -96 
NF protocol training | -96 
NF protocol awareness | -96 
NF protocol empowerment | -96 
NF protocol support | -96 
NF guideline safety | -96 
NF guideline education | -96 
NF guideline training | -96 
NF guideline awareness | -96 
NF guideline empowerment | -96 
NF guideline support | -96 
NF algorithm safety | -96 
NF algorithm education | -96 
NF algorithm training | -96 
NF algorithm awareness | -96 
NF algorithm empowerment | -96 
NF algorithm support | -96 
NF decision-making safety | -96 
NF decision-making education | -96 
NF decision-making training | -96 
NF decision-making awareness | -96 
NF decision-making empowerment | -96 
NF decision-making support | -96 
NF communication safety | -96 
NF communication education | -96 
NF communication training | -96 
NF communication awareness | -96 
NF communication empowerment | -96 
NF communication support | -96 
NF teamwork safety | -96 
NF teamwork education | -96 
NF teamwork training | -96 
NF teamwork awareness | -96 
NF teamwork empowerment | -96 
NF teamwork support | -96 
NF handoff safety | -96 
NF handoff education | -96 
NF handoff training | -96 
NF handoff awareness | -96 
NF handoff empowerment | -96 
NF handoff support | -96 
NF transition safety | -96 
NF transition education | -96 
NF transition training | -96 
NF transition awareness | -96 
NF transition empowerment | -96 
NF transition support | -96 
NF discharge safety | -96 
NF discharge education | -96 
NF discharge training | -96 
NF discharge awareness | -96 
NF discharge empowerment | -96 
NF discharge support | -96 
NF readmission safety | -96 
NF readmission education | -96 
NF readmission training | -96 
NF readmission awareness | -96 
NF readmission empowerment | -96 
NF readmission support | -96 
NF hospital-acquired condition | -96 
NF hospital-acquired infection | -96 
NF central line-associated bloodstream infection | -96 
NF catheter-associated urinary tract infection | -96 
NF ventilator-associated pneumonia | -96 
NF surgical site infection | -96 
NF pressure ulcer | -96 
NF fall | -96 
NF medication error | -96 
NF adverse drug reaction | -96 
NF allergic reaction | -96 
NF anaphylaxis | -96 
NF sentinel event | -96 
NF near miss | -96 
NF adverse event | -96 
NF root cause analysis | -96 
NF quality improvement initiative | -96 
NF patient safety initiative | -96 
NF patient safety goal | -96 
NF patient safety objective | -96 
NF patient safety target | -96 
NF patient safety metric | -96 
NF patient safety measure | -96 
NF patient safety benchmark | -96 
NF patient safety best practice | -96 
NF patient safety guideline | -96 
NF patient safety protocol | -96 
NF patient safety algorithm | -96 
NF patient safety decision-making | -96 
NF patient safety education | -96 
NF patient safety training | -96 
NF patient safety awareness | -96 
NF patient safety empowerment | -96 
NF patient safety support | -96 
NF family safety | -96 
NF family education | -96 
NF family training | -96 
NF family awareness | -96 
NF family empowerment | -96 
NF family support | -96 
NF healthcare provider safety | -96 
NF healthcare provider education | -96 
NF healthcare provider training | -96 
NF healthcare provider awareness | -96 
NF healthcare provider empowerment | -96 
NF healthcare provider support | -96 
NF staff safety | -96 
NF staff education | -96 
NF staff training | -96 
NF staff awareness | -96 
NF staff empowerment | -96 
NF staff support | -96 
NF leadership safety | -96 
NF leadership education | -96 
NF leadership training | -96 
NF leadership awareness | -96 
NF leadership empowerment | -96 
NF leadership support | -96 
NF management safety | -96 
NF management education | -96 
NF management training | -96 
NF management awareness | -96 
NF management empowerment | -96 
NF management support | -96 
NF governance safety | -96 
NF governance education | -96 
NF governance training | -96 
NF governance awareness | -96 
NF governance empowerment | -96 
NF governance support | -96 
NF policy safety | -96 
NF policy education | -96 
NF policy training | -96 
NF policy awareness | -96 
NF policy empowerment | -96 
NF policy support | -96 
NF procedure safety | -96 
NF procedure education | -96 
NF procedure training | -96 
NF procedure awareness | -96 
NF procedure empowerment | -96 
NF procedure support | -96 
NF protocol safety | -96 
NF protocol education | -96 
NF protocol training | -96 
NF protocol awareness | -96 
NF protocol empowerment | -96 
NF protocol support | -96 
NF guideline safety | -96 
NF guideline education | -96 
NF guideline training | -96 
NF guideline awareness | -96 
NF guideline empowerment | -96 
NF guideline support | -96 
NF algorithm safety | -96 
NF algorithm education | -96 
NF algorithm training | -96 
NF algorithm awareness | -96 
NF algorithm empowerment | -96 
NF algorithm support | -96 
NF decision-making safety | -96 
NF decision-making education | -96 
NF decision-making training | -96 
NF decision-making awareness | -96 
NF decision-making empowerment | -96 
NF decision-making support | -96 
NF communication safety | -96 
NF communication education | -96 
NF communication training | -96 
NF communication awareness | -96 
NF communication empowerment | -96 
NF communication support | -96 
NF teamwork safety | -96 
NF teamwork education | -96 
NF teamwork training | -96 
NF teamwork awareness | -96 
NF teamwork empowerment | -96 
NF teamwork support | -96 
NF handoff safety | -96 
NF handoff education | -96 
NF handoff training | -96 
NF handoff awareness | -96 
NF handoff empowerment | -96 
NF handoff support | -96 
NF transition safety | -96 
NF transition education | -96 
NF transition training | -96 
NF transition awareness | -96 
NF transition empowerment | -96 
NF transition support | -96 
NF discharge safety | -96 
NF discharge education | -96 
NF discharge training | -96 
NF discharge awareness | -96 
NF discharge empowerment | -96 
NF discharge support | -96 
NF readmission safety | -96 
NF readmission education | -96 
NF readmission training | -96 
NF readmission awareness | -96 
NF readmission empowerment | -96 
NF readmission support | -96 
NF hospital-acquired condition | -96 
NF hospital-acquired infection | -96 
NF central line-associated bloodstream infection | -96 
NF catheter-associated urinary tract infection | -96 
NF ventilator-associated pneumonia | -96 
NF surgical site infection | -96 
NF pressure ulcer | -96 
NF fall | -96 
NF medication error | -96 
NF adverse drug reaction | -96 
NF allergic reaction | -96 
NF anaphylaxis | -96 
NF sentinel event | -96 
NF near miss | -96 
NF adverse event | -96 
NF root cause analysis | -96 
NF quality improvement initiative | -96 
NF patient safety initiative | -96 
NF patient safety goal | -96 
NF patient safety objective | -96 
NF patient safety target | -96 
NF patient safety metric | -96 
NF patient safety measure | -96 
NF patient safety benchmark | -96 
NF patient safety best practice | -96 
NF patient safety guideline | -96 
NF patient safety protocol | -96 
NF patient safety algorithm | -96 
NF patient safety decision-making | -96 
NF patient safety education | -96 
NF patient safety training | -96 
NF patient safety awareness | -96 
NF patient safety empowerment | -96 
NF patient safety support | -96 
NF family safety | -96 
NF family education | -96 
NF family training | -96 
NF family awareness | -96 
NF family empowerment | -96 
NF family support | -96 
NF healthcare provider safety | -96 
NF healthcare provider education | -96 
NF healthcare provider training | -96 
NF healthcare provider awareness | -96 
NF healthcare provider empowerment | -96 
NF healthcare provider support | -96 
NF staff safety | -96 
NF staff education | -96 
NF staff training | -96 
NF staff awareness | -96 
NF staff empowerment | -96 
NF staff support | -96 
NF leadership safety | -96 
NF leadership education | -96 
NF leadership training | -96 
NF leadership awareness | -96 
NF leadership empowerment | -96 
NF leadership support | -96 
NF management safety | -96 
NF management education | -96 
NF management training | -96 
NF management awareness | -96 
NF management empowerment | -96 
NF management support | -96 
NF governance safety | -96 
NF governance education | -96 
NF governance training | -96 
NF governance awareness | -96 
NF governance empowerment | -96 
NF governance support | -96 
NF policy safety | -96 
NF policy education | -96 
NF policy training | -96 
NF policy awareness | -96 
NF policy empowerment | -96 
NF policy support | -96 
NF procedure safety | -96 
NF procedure education | -96 
NF procedure training | -96 
NF procedure awareness | -96 
NF procedure empowerment | -96 
NF procedure support | -96 
NF protocol safety | -96 
NF protocol education | -96 
NF protocol training | -96 
NF protocol awareness | -96 
NF protocol empowerment | -96 
NF protocol support | -96 
NF guideline safety | -96 
NF guideline education | -96 
NF guideline training | -96 
NF guideline awareness | -96 
NF guideline empowerment | -96 
NF guideline support | -96 
NF algorithm safety | -96 
NF algorithm education | -96 
NF algorithm training | -96 
NF algorithm awareness | -96 
NF algorithm empowerment | -96 
NF algorithm support | -96 
NF decision-making safety | -96 
NF decision-making education | -96 
NF decision-making training | -96 
NF decision-making awareness | -96 
NF decision-making empowerment | -96 
NF decision-making support | -96 
NF communication safety | -96 
NF communication education | -96 
NF communication training | -96 
NF communication awareness | -96 
NF communication empowerment | -96 
NF communication support | -96 
NF teamwork safety | -96 
NF teamwork education | -96 
NF teamwork training | -96 
NF teamwork awareness | -96 
NF teamwork empowerment | -96 
NF teamwork support | -96 
NF handoff safety | -96 
NF handoff education | -96 
NF handoff training | -96 
NF handoff awareness | -96 
NF handoff empowerment | -96 
NF handoff support | -96 
NF transition safety | -96 
NF transition education | -96 
NF transition training | -96 
NF transition awareness | -96 
NF transition empowerment | -96 
NF transition support | -96 
NF discharge safety | -96 
NF discharge education | -96 
NF discharge training | -96 
NF discharge awareness | -96 
