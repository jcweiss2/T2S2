67 years old | 0
male | 0
neck pain | -2160
ground-level fall | -2160
no signs or symptoms of radiculopathy | -2160
no signs or symptoms of myelopathy | -2160
5/5 strength on manual motor testing | -2160
normal sensation to light touch at the occiput | -2160
decreased sensation to light touch involving the right ear, face, and neck | -2160
normal upper and lower extremity reflexes | -2160
negative Hoffman’s sign | -2160
negative plantar Babinski reflex | -2160
negative Romberg sign | -2160
normal tandem gait | -2160
radiographs of the cervical spine | -2160
no evidence of pathology involving the cervical spine | -2160
persistent neck pain | -2160
CT scan of the cervical spine | -2160
destructive lesion with peripheral sclerosis involving the C2 body and odontoid | -2160
destruction of the posterior wall of the vertebral body | -2160
magnetic resonance imaging scan of the cervical spine | -2160
T2 hyperintense enhancing mass centered in the C2 body | -2160
extradural extension that displaced the spinal cord | -2160
no evidence of myelomalacia | -2160
mass extended into the odontoid, anterior arch and right lateral mass of C1, right C2–3 neural foramen, and right transverse process of C3 | -2160
complete encasement of the right vertebral artery | -2160
chordoma diagnosis | -2160
CT-guided needle biopsy | -2160
pathology review of the tissue specimen consistent with chordoma | -2160
CT scan of the chest, abdomen, and pelvis | -2160
no evidence of metastatic disease | -2160
en bloc tumor excision | 0
circumferential fusion | 0
reconstruction of the anterior column with free vascularized fibular grafting | 0
temporary balloon occlusion of the right vertebral artery | 0
embolization of the right vertebral artery | 0
surgery | 0
prone position | 0
Mayfield head holder | 0
corticocancellous struts and cancellous autograft from the right iliac crest | 0
exposure of the spine | 0
plane developed within the paraspinal muscles | 0
ligation of the right vertebral artery | 0
complete laminectomy at C1 | 0
partial laminectomies at C2 and C3 | 0
osteotomies through the lateral mass of C2 and the vertebral body of C3 | 0
transection of the right C2 and C3 nerve roots | 0
posterior instrumentation | 0
occipital plate | 0
3.5-mm screws bilaterally at C4 through C7 | 0
3.5-mm cobalt chrome rods bilaterally | 0
rib allograft and fibular allograft struts | 0
cancellous iliac crest autograft | 0
iliac crest strut graft | 0
postoperative care in the ICU | 0
disoriented | 24
unable to follow commands | 24
moving all 4 extremities sluggishly | 24
CT scan of the head | 24
new high-attenuation material within bilateral cerebellar hemispheres | 24
remote cerebellar hemorrhage | 24
interval repeat CT scans of the head | 48
no increase in the degree of hemorrhage | 48
progressive recovery of neurological function | 48
febrile | 120
worsening leukocytosis | 120
global decline in strength and mentation | 120
surgical incisions appeared benign | 120
CT scan of the neck with contrast | 120
right-sided anterior and posterior fluid collections | 120
concern for possible seromas, abscesses, or cerebrospinal fluid collections | 120
aspiration of fluid collections | 120
ultrasound-guided drains | 120
fluid from the drains returned positive for beta-2 transferrin | 120
bacterial cultures grew multiple colonies of Serratia marcescens | 120
inaccessible dural tear | 120
decision to remove the drains | 120
oversew the drain sites in a water-tight fashion | 120
lifelong antibiotic suppression | 120
severe dysphagia | 120
nasogastric tube feeds | 120
percutaneous endoscopic gastrostomy tube | 600
tracheostomy decannulation | 600
discharged home from the rehabilitation unit | 768
post-hospitalization course | 768
CT scan at 3 months postoperatively | 936
evidence of early osseous bridging | 936
severe dysphagia | 936
complete inability to tolerate food or liquid by mouth | 936
lifelong suppressive antibiotics | 936
physical examination | 936
intact strength in all key motor groups | 936
CT scan at 5 months postoperatively | 1200
complete fusion of the FVFG to the clivus and C4 | 1200
continued interval healing of the posterior strut grafts | 1200
no evidence of hardware failure | 1200
halo vest removal | 1200
isometric neck exercises | 1200
proton beam radiation | 1296
interval follow-up | 1296
no evidence of tumor recurrence | 1296
solid circumferential arthrodesis | 1296
follow-up endoscopic swallow evaluation | 4032
concern for thinning of the posterior pharyngeal wall | 4032
plate removal | 4032
repeat endoscopy | 4224
significant improvement in the gross appearance of the posterior pharyngeal wall | 4224
Neck Disability Index improvement | 8760
death from an unrelated medical condition | 10512