47 years old | 0
female | 0
admitted to the oncology ward | 0
low abdominal pain | -720
nausea | -720
vomiting | -720
hyporexia | -720
dehydration | -720
weight loss | -720
hypogastric mass | 0
ascites | 0
deep venous thrombosis (DVT) | 0
asymmetric edema | 0
anemia | 0
normal electrolytes | 0
preserved renal function | 0
preserved hepatic function | 0
pelvic mass | 0
infiltrating the left hepatic lobe | 0
peritoneum involvement | 0
multiple para-aortic and iliac lymph nodes | 0
bilateral pleural effusion | 0
neoplastic cells in pleural and ascitic fluids | 0
image-guided biopsy of a peritoneal nodule | 0
poorly differentiated small-cell neoplasia | 0
immunohistochemistry analysis | 0
positive for CD56 | 0
positive for vimentin | 0
focally positive for cytokeratins 35BH11 | 0
negative for WT1 | 0
negative for estrogen receptor | 0
negative for TTF-1 | 0
negative for inhibin | 0
carcinoma with neuroendocrine differentiation | 0
ovarian biopsy | 28
emergency laparotomy | 28
acute peritonitis | 28
septic shock | 35
febrile neutropenia | 35
necrotic adnexal mass | 35
abscess | 35
venous hydration | 0
anticoagulation with low-molecular weight heparin | 0
systemic chemotherapy | 0
cisplatin | 0
etoposide | 0
remarkable clinical response | 21
reduction of the abdominal mass | 21
improvement of performance status | 21
tumor lysis syndrome (TLS) | 2
hyperkalemia | 2
hyperphosphatemia | 2
hypocalcemia | 2
second chemotherapy cycle | 28
sepsis | 35
death | 42