11 years old | 0
girl | 0
admitted to the hospital | 0
fever | -72
vomiting | -72
generalized abdominal pain | -72
rash on palms | 0
rash on trunk | 0
severe drowsiness | 0
lethargic | 0
no conjunctivitis | 0
no lymphadenopathy | 0
respiratory rate 25/min | 0
oxygen saturation 93% | 0
harsh breathing with crackles during inspiration | 0
tachycardia (HR 135 bpm) | 0
hypotension (BP 80/42 mm Hg) | 0
abdomen tender to palpation (right lower quadrant) | 0
white blood cell count 13.5 ×103/μL | 0
neutrophils 94.5% | 0
erythrocyte sedimentation rate 82 mm/h | 0
CRP 298.5 mg/L | 0
procalcitonin 18.45 mcg/L | 0
negative SARS-CoV-2 PCR | 0
negative SARS-CoV-2 RT-PCR | 0
abdominal ultrasound enlarged appendix (11.2 mm) | 0
fluid in pelvis | 0
emergency laparotomy appendectomy | 0
postoperative tachycardia (139 bpm) | 0
postoperative hypotension (BP 76/39 mmHg) | 0
fractional shortening on echocardiogram | 0
oxygen saturation 88-90% | 0
oxygen therapy (2 L/min O2) | 0
chest X-ray bilateral paratracheal and paracardial spots | 0
ceftriaxone treatment | 0
amikacin treatment | 0
imipenem treatment | 0
history of contact with COVID-19 (grandfather) | -720
positive SARS-CoV-2 IgG | 24
elevated ferritin | 24
elevated IL6 | 24
elevated high-sensitivity troponin | 24
elevated D-dimer | 24
enoxaparin treatment | 24
IVIG treatment | 24
aspirin treatment | 24
hemoglobin decreased (11.5 to 6.9 g/dL) | 48
red blood cell transfusion | 48
methylprednisolone treatment | 48
LV dysfunction (EF 30%) | 48
dobutamine treatment | 48
afebrile | 96
arterial pressure stable | 96
no pathogenic agents detected in cultures | 96
catarrhal appendicitis diagnosis | 96
D-dimer downward trend | 96
troponemia resolved | 96
inflammatory parameters normal | 96
LV function improved | 96
discharge | 288
low-dose aspirin (3 mg/kg) | 288
blood tests normalized | 336
COV-2 IgG elevated (84) | 336
abdominal ultrasound normal | 336
cardiac ultrasound normal | 336
follow-up every 3 months | 336
no short-term complications | 336
