50 years old | 0
male | 0
admitted to the hospital | 0
edema of the legs | 0
erythema | 0
pain | 0
abdominal swelling | 0
pulmonary hypertension | 0
right heart failure | 0
atrial fibrillation | 0
chronic obstructive pulmonary disease | 0
cellulitis | 0
history of appendectomy | -10800
stabbed in the abdomen | -5400
treated by general surgery | -5400
discharged from hospital | -5393
history of smoking | -14400
shortness of breath | -1800
diagnosed with NYHA Class II | -1800
echocardiography | -1800
right heart cavity dimensions mildly increased | -1800
pulmonary artery systolic pressure 45 mmHg | -1800
treated and complaints regressed | -1800
admitted to the Pulmonology department | -1080
abdominal and bilateral leg swelling | -1080
shortness of breath | -1080
diagnosed with right heart failure | -1080
CT thorax | -1080
treated with diuretics, steroids, theophylline, and inhaled bronchodilator | -1080
complaints regressed | -1080
echo findings | -1080
left ventricular ejection fraction 65% | -1080
Grade I diastolic dysfunction | -1080
normal left heart cavities | -1080
significantly enlarged right heart cavities | -1080
pulmonary artery systolic pressure 70 mmHg | -1080
Grade 2-3 tricuspid failure | -1080
admitted to the Pulmonology department | -720
high ventricular rate atrial fibrillation | -720
abdominal ascites | -720
diffuse edema of the lower extremities | -720
crackles in the middle and lower lung zones | -720
NYHA functional Class IV | -720
treated with digoxin, diltiazem, and warfarin | -720
symptoms regressed to NYHA Class III | -720
discharged from hospital | -713
admitted to Emergency department | -695
worsening right heart failure | -695
shortness of breath | -695
transferred to the Cardiology department | -695
treated with intravenous furosemide, spironolactone, clexane, diltiazem, and digoxin | -695
started on ampicillin/sulbactam | -695
laboratory findings | -695
blood urea nitrogen 60 mg/dl | -695
creatinine 1.2 mg/dl | -695
aspartate aminotransferase 40 U/l | -695
alanine aminotransferase 45 U/l | -695
hemoglobin 12.8 g/dl | -695
white blood cells 14,500/µl | -695
respiratory arrest | 48
cardiac arrest | 48
cardiopulmonary resuscitation | 48
intubated | 48
basal rhythm of atrial fibrillation | 48
blood pressure 100/60 mmHg | 48
transferred to the intensive care unit | 48
mechanic ventilator | 48
pulmonary CT angiography | 48
no thrombi detected | 48
CT thorax angiography | 48
lower extremity venous Doppler ultrasonography | 48
no thrombotic formation detected | 48
abdominal auscultation | 48
diagnosis of aortocaval fistula | 48
IVC diameter 19 cm | 48
harsh pansystolic murmur | 48
liver palpable 7-8 cm under the costal arch | 48
diffuse ascites | 48
edema of the legs 3+ | 48
continuous thrill and machine-like murmur | 48
echo findings | 48
right cardiac cavities severely enlarged | 48
3-4 degree of tricuspid failure | 48
pulmonary artery pressure 75-80 mmHg | 48
normal left heart cavities | 48
IVC measured 18 cm | 48
fistula between the abdominal aorta and the IVC | 48
transesophageal echocardiography | 48
intact interventricular septum | 48
patent foramen ovale | 48
right to left shunt | 48
CT angiography | 48
fistula between the abdominal aorta and the IVC | 48
diameter of the aorta 22 mm | 48
IVC diameter 99 mm | 48
diameter of the fistula tract 11 mm | 48
diameter of the aorta 25 mm | 48
IVC diameter 169 mm | 48
fistula tract diameter 17 mm | 48
abdominal aortography | 48
findings consistent with CT angiography | 48
oxymetrically calculated left-to-right shunt 2.8 | 48
coronary angiography | 48
coronary arteries normal | 48
systolic pulmonary artery pressure 75 mmHg | 48
decision to close the ACP percutaneously | 48
pneumonia did not resolve | 120
developed sepsis | 120
died of septic shock | 120