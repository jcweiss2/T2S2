27 years old | 0
female | 0
Gravida 4 | 0
Para 3 | 0
17 weeks gestation | 0
admitted to the hospital | 0
fever | -72
dry cough | -72
shortness of breath | -72
diagnosed with COVID-19 | -72
COVID-19 vaccine dose | -264
body temperature 39.0 °C | 0
oxygen saturation 84% | 0
respiratory rate 30 breaths/minute | 0
blood pressure 130/80 mmHg | 0
pulse 125 beats per minute | 0
transferred to ICU | 0
high-flow nasal cannula | 0
fraction of inspired oxygen 100% | 0
bilevel positive airway pressure | 24
expiratory positive airway pressure 8 cmH2O | 24
inspiratory positive airway pressure 13 cmH2O | 24
intubated | 96
invasive mechanical ventilation | 96
dexamethasone 6 mg/day | 0
enoxaparin 60 mg twice a day | 0
clopidogrel 75 mg daily | 0
ceftriaxone 2 g/day | 0
multivitamin | 0
magnesium | 0
zinc | 0
nasal gastric enteral feeding | 0
parenteral nutrition | 0
therapeutic plasma exchange | 144
human albumin replacement | 144
improved clinical status | 168
improved arterial blood gas | 168
improved biochemical parameters | 168
fever 39 °C | 288
antibiotic treatment changed | 288
extubated | 312
CPAP | 312
fraction of inspired oxygen 60% | 312
high-flow nasal cannula | 360
fraction of inspired oxygen 33% | 360
oxygen support discontinued | 504
discharged from hospital | 648
healthy 20-week gestational fetus | 648