7 days old | 0
female | 0
admitted to the hospital | 0
poor feeding | -24
bloody stools | -24
loss of consciousness | -18
transported to NICU | -18
temperature 35.6°C | 0
heart rate 170 beats per minute | 0
respiratory rate 65 times per minute | 0
capillary refill time >3 seconds | 0
blood pressure 35/23mmHg | 0
unresponsive | 0
dry mucous membranes |,0
diminished pulses | 0
mottled cold extremities | 0
decreased urine output | 0
significant abdominal distention | 0
WBC 38.51×109/L | 0
polymorphonuclear cells 49% | 0
lymphocytes 38.8% | 0
monocytes 12.2% | 0
hemoglobin 14.6g/dL | 0
platelet count 279×109/L | 0
C-reactive protein 37mg/L | 0
prothrombin time 16.2 sec | 0
activated partial thromboplastin time 34 sec | 0
necrotizing enterocolitis | 0
pneumatosis intestinalis | 0
portal venous gas | 0
ascitic fluid WBC count 2815×106/L | 6
ascitic fluid polymorphonuclear cells 56% | 6
ascitic fluid lymphocytes 15% | 6
ascitic fluid monocytes/macrophages 29% | 6
ascitic fluid red blood cell count 55×106/L | 6
blood culture no bacterial growth | 0
fecal culture no bacterial growth | 0
normal saline administration | 0
dopamine administration | 0
ceftazidime | 0
penicillin G sodium | 0
abdominal distension increased | 2
soy sauce-colored urine | 2
jaundice | 2
hemoglobin decrease 14.6 g/dL to 5.1 g/dL | 2
direct antiglobulin test negative | 2
acid elution negative | 2
red blood cell transfusion | 2
blood potassium 8.7mmol/L | 2
premature ventricular contractions | 2
continuous renal replacement therapy | 2
vancomycin | 2
meropenem | 2
prothrombin time >180 sec | 11
activated partial thromboplastin time >120 sec | 11
fibrin degradation products increase | 11
D-Dimer increase | 11
disseminated intravascular coagulation | 11
metagenomic next-generation sequencing positive for C. perfringens | 18
multi-organ failure | 18
death | 48
