79 years old | 0
male | 0
hypertension | 0
ischemic heart disease | 0
admitted to the hospital | 0
severe symptomatic aortic stenosis | 0
coronary artery bypass graft surgery | -132
mitral valve repair | -132
preprocedural transthoracic echocardiography | -1
severe aortic stenosis | -1
left ventricular ejection fraction of 45% | -1
induction of general anesthesia | 0
TEE probe insertion | 0
SAPIEN 3 valve deployment | 0
postprocedural TEE | 1
prosthesis in good position | 1
no visible paravalvular leak | 1
gastric aspiration with an orogastric tube | 1
blood-tinged secretions | 1
extubated | 1
transferred to the intensive care unit | 1
progressive chest pain | 2
important shivering | 2
computed tomography (CT) with intravenous contrast | 2
pneumomediastinum | 2
right hydropneumothorax | 2
esophageal perforation suspected | 2
right thoracic drain inserted | 2
serosanguinous liquid drained | 2
esophagogastroscopy | 2
4-cm vertical perforation of the middle third of the esophagus | 2
returned to the operating room | 7
right thoracotomy | 7
repair of an esophageal perforation | 7
lysis of extensive pleural adhesions | 7
esophageal laceration site found | 7
large vertebral osteophyte visualized | 7
primary closure of the esophageal wall | 7
intercostal muscular flap mobilized | 7
thoracic drains left in place | 7
transferred to the intensive care unit | 7
pneumonia | 24
severe delirium | 24
congestive heart failure with pulmonary edema | 24
died after withdrawal of care | 720