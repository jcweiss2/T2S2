58 years old | 0
male | 0
schizophrenia | 0
substance abuse | 0
diabetes mellitus | 0
hypertension | 0
admitted to the hospital | 0
headache | 0
chest pain | 0
afebrile | 0
hypertensive | 0
tachycardic | 0
confused | 0
intubated | 0
hyperglycemia | 0
acute kidney injury | 0
creatinine 1.6 | 0
baseline creatinine 1.1 | 0
extubated | 24
altered mental status attributed to synthetic cannabinoid intoxication | 24
increasingly agitated | 96
tachycardic | 96
hypertensive | 96
abdominal distension increased | 96
progressively hypotensive | 144
intravenous fluid resuscitation | 144
febrile | 192
re-intubated | 192
respiratory distress | 192
arterial lactate peaked at 2.1 mmol/L | 192
empirically treated with piperacillin-tazobactam | 192
blood cultures grew Lactobacillus species | 192
persistent bandemia | 192
worsening diarrhea | 192
metronidazole added | 192
noncontrast CT showed wall thickening of the ascending colon | 192
ileus | 192
C. difficile toxin in stool negative | 192
colonoscopy showed diffuse edema | 192
severe ulceration | 192
necrotic mucosa | 192
ischemic colitis | 192
transesophageal echocardiogram showed no vegetation | 192
improved clinically | 336
extubated | 336
discharged | 336