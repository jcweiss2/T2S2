27 years old | 0
male | 0
admitted to the emergency department | 0
diffuse abdominal pain | -24
multiple episodes of vomiting of gastric content | -24
blunt abdominal trauma caused by a kick with a knee to the abdomen | -24
high heart rate of 94 beats/min | 0
respiratory rate of 19 breaths/min | 0
blood pressure of 130/50 mmHg | 0
temperature 36 °C | 0
oxygen saturation level of 94 % | 0
generalized abdominal pain on palpation | 0
predominant pain in the lower abdomen | 0
voluntary muscular defense | 0
signs of peritoneal irritation | 0
normal hemoglobin level | 0
mild leukocytosis | 0
hemoglobin: 17.6 g/dL | 0
hematocrit: 52 % | 0
leukocytes: 13.1 × 10³/μL | 0
platelets: 317 × 10³/μL | 0
creatinine within normal limits | 0
urinalysis within normal limits | 0
computed tomography showing rupture of the third portion of the duodenum | 0
computed tomography showing retropneumoperitoneum | 0
exploratory laparotomy | 0
free perforation of approximately 1 cm in the posterior wall of the third portion of the duodenum | 0
Kocher maneuver | 0
duodenorrhaphy with Connel-Mayo suture | 0
Lambert suture with vascular prolene | 0
Jackson-Pratt drain placement | 0
nasogastric tube placement | 0
peritoneal fluid culture | 0
Gram stain of peritoneal fluid | 0
piperacillin-tazobactam antibiotic coverage | 0
enteral nutrition for one week | 168
drain removal | 360
peritoneal fluid culture reported Enterobacter cloacae complex | 168
inducible strain producing beta-lactamases | 168
AmpC pattern | 168
evaluation by infectology service | 168
ertapenem titration over 10 days | 168
elevated acute phase reactants | 168
leukocytosis | 168
postoperative control a week later | 168
postoperative control one month later | 672
early diet recommendation | 168
physical therapy recommendation | 168
early mobilization recommendation | 168
restricted sports activity for one month | 672
hospitalized for three weeks | 504
secondary peritonitis | 0
uncontained perforation | 0
pneumoperitoneum | 0
free perforation | 0
contamination in peritoneal cavity | 0
closure of duodenal lesion | 0
discharge | 504
