60 years old | 0
female | 0
abdominal incisional hernia | -5 years
laparotomic appendectomy | -5 years
acute appendicitis | -5 years
peritoneal abscess | -5 years
abdominal wall bulging | 0
xipho-pubic scar | 0
tumefaction | 0
abdominoplasty | 0
incisional hernia repair | 0
open keel technique | 0
xipho-pubic scar excised | 0
dissection of the umbilicus | 0
supra-umbilical hernia sac dissection | 0
linear median incision | 0
viscerolysis | 0
abdominal wall defect correction | 0
rectus abdominis muscle plasty | 0
umbilicus reconstruction | 0
Redon type surgical drains placement | 0
weak peristalsis | 48
afebrile | 48
good general conditions | 48
deambulation | 48
bowels open | 72
drains removed | 96
discharged | 96
follow-up | 100
clean healing wound | 100
deterged and dressed | 100
stitches removed | 552
median epigastric bulge | 696
fever | 696
ballottement | 696
erythema | 696
pain | 696
pus drained | 696
subcutaneous abscess | 696
antibiotic therapy | 698
persistent pain | 744
xipho-umbilical bulge | 744
purulent exudate | 744
dyspnoea | 744
chest X-ray | 744
abdominal CT scan | 744
intestinal perforation | 744
exploratory laparotomy | 744
plastic peritonitis | 744
extended right and transverse colectomy | 744
perforation and abscessing mass | 744
right monolateral salpingo-ovariectomy | 744
temporary ileostomy | 744
histological examination | 744
haemorrhagic serositis | 744
ischaemic necrosis | 744
ulceration | 744
postoperative care | 744
Metronidazole administration | 744
Levofloxacin administration | 744
Imipenem administration | 744
Tigecicline administration | 744
Fluconazole administration | 744
ileostomy reversal surgery | 900
discharged | 944