57 years old | 0
female | 0
presented to the emergency department | -72
acute abdominal pain | -72
acute in onset | -72
crampy pain | -72
non-radiating pain | -72
pain increasing in severity | -72
pain aggravated after ingestion of food | -72
palpitation | -72
vomiting | -72
vomiting episodes | -48
no stool passage | -48
no flatus passage | -48
chronic smoker | -87600
Chronic Obstructive Pulmonary Disease | -87600
pulse rate 130 beats per minute | 0
regular pulse | 0
oxygen saturation 85% on room air | 0
blood pressure 95/70 mm Hg | 0
body temperature 38.7 °C | 0
respiratory rate 22 breaths/min | 0
sinus rhythm tachycardia | 0
rapid antigen test positive | 0
RT-PCR positive | 0
distended abdomen | 0
diffuse tenderness | 0
diffuse guarding | 0
rigidity | 0
absent bowel sounds | 0
normal sphincter tone | 0
collapsed rectum | 0
absent fecal stain | 0
crystalloids administered | 0
supplemental oxygen 4 L/min | 0
nasogastric tube decompression | 0
Foley catheterization | 0
leukocytosis | 0
raised amylase | 0
total bilirubin 2.20 mg/dL | 0
conjugated bilirubin 0.9 mg/dL | 0
alkaline phosphatase 674 U/L | 0
metabolic acidosis | 0
raised lactate level | 0
WBC count 13 ×10^9 cells/L | 0
neutrophil 80% | 0
lymphocyte 15% | 0
hemoglobin 13.3 g/dL | 0
platelet count 229 ×10^9 cells/L | 0
total bilirubin 2.2 mg/dL | 0
direct bilirubin 0.9 mg/dL | 0
AST 10 U/L | 0
ALT 15 U/L | 0
albumin 3.9 g/L | 0
amylase 216 U/L | 0
lipase 58 U/L | 0
blood sodium 138 mEq/L | 0
blood potassium 4.4 mEq/L | 0
blood calcium 6.9 mg/dL | 0
blood urea nitrogen 54 mg/dL | 0
creatinine 0.6 mg/dL | 0
FDP D-dimer 0.8 μg/mL | 0
prominent dilated small bowel loops | 0
absence of completely visible colon | 0
multiple air fluid levels | 0
small bowel obstruction | 0
minimal free fluid in pelvis | 0
fluid collection in right iliac fossa | 0
fluid collection in pelvis | 0
fluid collection along anterior liver surface | 0
emergency laparotomy | 0
greenish fluid | 0
gangrenous small bowel | 0
tissue decay | 0
blackish discoloration of intestine | 0
AMI | 0
resection of gangrenous bowel | 0
double barrel loop ileostomy | 0
shifted to COVID ICU | 0
Meropenem IV 1 g | 24
Vancomycin IV 500 mg | 24
low molecular weight Heparin 60 mg | 24
total parenteral nutrition | 24
small bowel necrosis | 24
microthrombi in lamina propria | 24
microthrombi in submucosa | 24
glandular necrosis | 24
COVID pneumonia | 144
reintubated | 144
sepsis | 144
Acute Kidney Injury | 144
expired | 336
severe sepsis | 336
multi-organ dysfunction syndrome | 336
57 years old|0
female|0
presented to the emergency department|-72
acute abdominal pain|-72
acute in onset|-72
crampy pain|-72
non-radiating pain|-72
pain increasing in severity|-72
pain aggravated after ingestion of food|-72
palpitation|-72
vomiting|-72
vomiting episodes|-48
no stool passage|-48
no flatus passage|-48
chronic smoker|-87600
Chronic Obstructive Pulmonary Disease|-87600
pulse rate 130 beats per minute|0
regular pulse|0
oxygen saturation 85% on room air|0
blood pressure 95/70 mm Hg|0
body temperature 38.7 °C|0
respiratory rate 22 breaths/min|0
sinus rhythm tachycardia|0
rapid antigen test positive|0
RT-PCR positive|0
distended abdomen|0
diffuse tenderness|0
diffuse guarding|0
rigidity|0
absent bowel sounds|0
normal sphincter tone|0
collapsed rectum|0
absent fecal stain|0
crystalloids administered|0
supplemental oxygen 4 L/min|0
nasogastric tube decompression|0
Foley catheterization|0
leukocytosis|0
raised amylase|0
total bilirubin 2.20 mg/dL|0
conjugated bilirubin 0.9 mg/dL|0
alkaline phosphatase 674 U/L|0
metabolic acidosis|0
raised lactate level|0
WBC count 13 ×10^9 cells/L|0
neutrophil 80%|0
lymphocyte 15%|0
hemoglobin 13.3 g/dL|0
platelet count 229 ×10^9 cells/L|0
total bilirubin 2.2 mg/dL|0
direct bilirubin 0.9 mg/dL|0
AST 10 U/L|0
ALT 15 U/L|0
albumin 3.9 g/L|0
amylase 216 U/L|0
lipase 58 U/L|0
blood sodium 138 mEq/L|0
blood potassium 4.4 mEq/L|0
blood calcium 6.9 mg/dL|0
blood urea nitrogen 54 mg/dL|0
creatinine 0.6 mg/dL|0
FDP D-dimer 0.8 μg/mL|0
prominent dilated small bowel loops|0
absence of completely visible colon|0
multiple air fluid levels|0
small bowel obstruction|0
minimal free fluid in pelvis|0
fluid collection in right iliac fossa|0
fluid collection in pelvis|0
fluid collection along anterior liver surface|0
emergency laparotomy|0
greenish fluid|0
gangrenous small bowel|0
tissue decay|0
blackish discoloration of intestine|0
AMI|0
resection of gangrenous bowel|0
double barrel loop ileostomy|0
shifted to COVID ICU|0
Meropenem IV 1 g|24
Vancomycin IV 500 mg|24
low molecular weight Heparin 60 mg|24
total parenteral nutrition|24
small bowel necrosis|24
microthrombi in lamina propria|24
microthrombi in submucosa|24
glandular necrosis|24
COVID pneumonia|144
reintubated|144
sepsis|144
Acute Kidney Injury|144
expired|336
severe sepsis|336
multi-organ dysfunction syndrome|336
