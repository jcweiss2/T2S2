36 years old | 0
male | 0
admitted to the hospital | 0
low-grade fever | -96
sore throat | -96
myalgia | -96
nausea | -96
injected pharynx | 0
thrombocytopenia | 0
platelet of 45,000/uL | 0
hemoglobin of 14.8 g/dL | 0
cell count of 8700 cells/uL | 0
neutrophil of 85% | 0
band form of 6% | 0
elevated creatinine of 2.1 mg/dL | 0
diagnosed with viral upper respiratory tract infection | 0
received 2 L of intravenous normal saline | 0
high fever of 39.2°C | 48
pleuritic chest pain | 48
low blood pressure of 80/50 mmHg | 48
transferred to Intensive care unit | 48
resuscitated with intravenous fluids | 48
blood cultures were obtained | 48
empirical antibiotics | 48
vancomycin | 48
piperacillin/tazobactam | 48
bilateral patchy and irregular parenchymal opacities | 48
right-sided pleural effusion | 48
multiple thick-walled cavitary and nodular opacities | 48
septic emboli | 48
blood cultures grew F. necrophorum | 72
antibiotic therapy was narrowed down to piperacillin/tazobactam | 72
responded well to intravenous fluids and antibiotics | 72
normalized blood pressure | 72
received 5 L of intravenous normal saline | 72
venous duplex ultrasonography | 72
thrombus in the left IJV | 72
diagnosed with Lemierre's syndrome | 72
pleural effusion was managed conservatively | 72
piperacillin/tazobactam was continued for 7 days | 168
discharged home | 168
4-week course of intravenous ertapenem | 168
recovered well from the infection | 336
no anticoagulation | 0