68 years old | 0
male | 0
from New Jersey | 0
immigrated from South Asia | -14760
lifestyle-controlled diabetes mellitus | -720
hyperlipidemia | -720
L4-L5 radiculopathy | -720
decompressive laminectomy | -720
herniation | -720
Aspirin | -720
non-smoker | 0
does not abuse alcohol or drugs | 0
BMI 24.2 | 0
fatigue | -72
dyspnea | -72
cough | -72
chills | -72
fever | -72
Tmax 101oF | -72
frank hematuria | -48
hypoxic | -48
SpO2 high 80s | -48
febrile | -48
tested positive for COVID-19 | -48
acute kidney injury | -48
hydroxychloroquine | 0
azithromycin | 0
progressive dyspnea | 24
hypoxia | 24
severe hypotension | 24
blood pressures documented as low as 60/40 | 24
intubated | 24
central access | 24
common femoral artery | 24
transitioned to the intensive care unit | 24
increasing pressure requirements | 120
persistent fevers | 120
Tmax 103.5oF | 120
hypotension | 120
cytokine storm | 120
Tocilizumab | 120
stabilized hemodynamically | 168
self-extubation | 168
supplemental oxygen | 168
high-flow nasal cannula | 168
weaned to room air | 240
discharged to inpatient rehabilitation | 240
negative COVID-19 test result | 240
asymptomatic deep venous thrombosis | 288
common femoral vein | 288
prophylactic heparin | 288
therapeutic Enoxaparin sodium | 288
acute pain in the right knee | 408
limited range of motion | 408
could not bear weight | 408
knee swollen | 408
knee painful | 408
ultrasound | 408
7 cm suprapatellar joint effusion | 408
low-grade fever | 408
Tmax 100.8oF | 408
warm | 408
erythematous knee | 408
knee arthrocentesis | 408
orthopedic surgery | 408
septic arthritis | 408
80cc of synovial fluid | 408
mild improvement in pain | 408
readmitted to the hospital | 432
blood pressure of 121/68 | 432
heart rate of 68 beats/min | 432
respiration rate of 20 respirations/min | 432
temperature of 98.4oF | 432
empiric antibiotics | 432
Vancomycin | 432
Zosyn | 432
high white blood cell count | 432
high lymphocytes | 432
low monocytes | 432
IL markers elevated | 432
microscopic review of the aspirate | 432
cloudy yellow synovial fluid | 432
neutrophilic predominance of 87% | 432
no crystals | 432
bacterial culture showed no growth | 432
intravenous antibiotics | 432
oral cephalexin | 432
Prednisone taper | 432
IL aseptic arthropathy | 432
transferred back to inpatient rehabilitation | 432
weakness | 432
poor endurance | 432
hospitalization for severe illness | 432
therapeutic Enoxaparin sodium | 432
oral Apixaban | 432
discharged home | 504