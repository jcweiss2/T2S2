31 years old | 0
male | 0
admitted to the hospital | 0
laparoscopic cholecystectomy | -672
CBD exploration | -672
T-tube placement | -672
follow-up visit | -672
cholangiogram | -672
T-tube removal | 0
severe abdominal pain | 0
tachycardia | 0
admission to the hospital | 0
abdominal ultrasound | 0
small fluid collection | 0
conservative management | 0
ERCP | 24
bile leak | 24
rupture at the point where the fistulous tract joined the abdominal wall | 24
contrast material leaking into the abdominal cavity | 24
endoscopic sphincterotomy | 24
biliary stent | 24
fever | 48
diaphoresis | 48
leucocytosis | 48
acute abdomen | 48
emergency laparoscopy | 48
severe generalized biliary-purulent peritonitis | 48
extensive lavage | 48
placement of abdominal drains | 48
rupture of the fistulous tract sutured | 48
hemodynamic instability | 48
bacteremia | 48
transfer to the ICU | 48
severe respiratory distress | 48
systemic inflammatory response syndrome | 48
septic shock | 48
ventilatory support | 48
multiple antibiotics | 48
vasoactive agents | 48
activated C protein | 48
culture of the peritoneal fluid | 48
multiresistant Pseudomonas aeruginosa | 48
discharged | 360
T-tube choledochotomy | -100 years
laparoscopic cholecystectomy | -20 years
cholecystectomy | -20 years
CBD exploration | -20 years
T-tube placement | -20 years
ERCP | -20 years
endoscopic sphincterotomy | -20 years
biliary stent | -20 years
transcystic exploration | -10 years
pneumatic dilatation | -10 years
choledochoscope | -10 years
transcystic stent | -10 years
guidewire | -10 years
postoperative ERCP | -10 years
primary closure of the CBD | -5 years
endobiliary stent | -5 years
bilioenteric reconstruction | -5 years
fistulogram | -5 years