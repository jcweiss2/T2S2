82 years old | 0
male | 0
Caucasian | 0
ECOG PS 0 | 0
hypertension | -8760
tobacco consumption | -8760
alcohol consumption | -8760
progressive growth of axillary and cervical lymph nodes | -720
biopsy | -720
MCC lymph node metastasis | -720
CK20+ | -720
CK7- | -720
TTF1- | -720
chromogranin+ | -720
synaptophysin+ | -720
staging PET 68-Ga DOTANOC | -672
supradiaphragmatic lymph node metastases | -672
pembrolizumab treatment start | 0
pembrolizumab 2 mg/kg q3w | 0
objective clinical response | 96
acute anorexia | 96
mental confusion | 96
obnubilation | 96
dehydration | 96
hyperglycemia | 96
acute kidney injury grade 3 | 96
hyponatremia | 96
hypercalcemia | 96
hyperphosphatemia | 96
ketonuria | 96
respiratory arrest | 96
bradycardia | 96
hypotension | 96
orotracheal intubation | 96
mechanic ventilation | 96
aminergic support | 96
mixed metabolic acidemia | 96
diabetic ketoacidosis diagnosis | 96
insulin therapy start | 96
corticosteroid therapy start | 120
discharged | 336
basal bolus insulin therapy | 4320
dysarthria | 4320
ataxia | 4320
admission to Oncology Ward | 4320
chest-abdomen-pelvis computed tomography | 4320
substantial partial response | 4320
axillary lymph node metastasis | 4320
brain and neural-axis magnetic resonance imaging | 4320
electromyography | 4320
mild axonal sensorimotor polyneuropathy | 4320
ANA ≥1/640 | 4320
lumbar puncture analysis | 4320
slight proteinorachia | 4320
absent pleocytosis | 4320
intrathecal antibody synthesis | 4320
mirror banding profile | 4320
systemic inflammation | 4320
immunofluorescence assay | 4320
fine granular IgG staining | 4320
methylprednisolone pulse therapy | 4464
neurologic deficits worsening | 4536
appendicular and axial ataxia | 4536
cerebellar dysarthria | 4536
dysphagia | 4536
methylprednisolone and intravenous immunoglobulin | 4536
nasogastric tube placement | 4536
gastric mucosa infiltration | 4536
biopsies | 4536
carcinoma CK20+ | 4536
NSE+ | 4536
CD56+ | 4536
chromogranin A+ | 4536
synaptophysin+ | 4536
CD117+ | 4536
MCC progression | 4536
palliative care start | 4536
death | 4608