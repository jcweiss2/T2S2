87 years old | 0
male | 0
admitted to the hospital | 0
coronary artery disease | -8760
TIA | -8760
hypertension | -8760
hyperlipidemia | -8760
osteoporosis | -8760
glaucoma | -8760
smoked | -525600
quit smoking | -525600
bitten by dog | -72
cellulitis | -72
ampicillin/sulbactam | -72
amoxicillin/clavulanate | -72
follow up | -72
erythema | -72
edema | -72
warmth | -72
hospitalization | -72
intravenous ampicillin/sulbactam | -72
vancomycin | -72
improvement | -24
discharged | -24
amoxicillin | -24
minocycline | -24
ankle pain | 0
loose bowel movements | 0
fever | 0
hypotension | 0
tachycardia | 0
tachypnea | 0
low oxygen saturation | 0
crackles | 0
systolic murmur | 0
flat JVP | 0
mild erythema | 0
eschar | 0
mild ankle warmth | 0
mild ankle edema | 0
leukocytosis | 0
neutrophils | 0
lymphocytes | 0
eosinophils | 0
elevated creatinine | 0
normal liver enzymes | 0
bilateral effusions | 0
lung infiltrates | 0
diagnosed with ankle sprain | 0
severe sepsis | 0
pneumonia | 0
acute kidney injury | 0
intravenous ertapenem | 0
intravenous vancomycin | 0
intravenous azithromycin | 0
oral metronidazole | 0
worsening tachypnea | 48
worsening hypoxia | 48
supplemental oxygen | 48
eosinophilia | 48
leukocytosis | 48
repeat chest film | 48
diffuse alveolar filling pattern | 48
acute respiratory distress syndrome | 48
computed tomography of the chest | 48
diffuse bilateral airspace disease | 48
ground glass attenuation | 48
bilateral pleural effusions | 48
intubated | 72
flexible fiberoptic bronchoscopy | 72
BAL | 72
transbronchial biopsies | 72
mechanical ventilation | 72
pneumothorax | 96
chest tube | 96
streptococcus parasanguinus | 96
Klebsiella | 96
C. difficile toxin | 96
urine legionella antigen | 96
coccidioides IgG | 96
coccidioides IgM | 96
ampicillin/sulbactam | 96
ciprofloxacin | 96
BAL sample | 120
nucleated cells | 120
neutrophils | 120
lymphocytes | 120
eosinophils | 120
transbronchial biopsies | 120
methylprednisolone | 120
leukocytosis | 144
eosinophilia | 144
defervesced | 144
improvement in gas exchange | 144
liberated from mechanical ventilation | 144
supplemental oxygen | 144
normalization of eosinophilia | 144
improvement in air space disease | 144
oral prednisone | 144
ciprofloxacin discontinued | 144
chest tube removed | 360
transthoracic echocardiogram | 360
no endocarditis | 360
sterile blood cultures | 360
vancomycin completed | 360
rehabilitation | 720
discharged | 720
follow up | 8760
no respiratory symptoms | 8760
inhaled mometasone | 8760
prednisone taper | 8760