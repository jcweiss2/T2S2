59 years old | 0
woman | 0
severe mitral valve insufficiency | 0
underwent MVR surgery | -87600
severe dysfunction of her prosthetic mitral valve | 0
redo MVR | 0
symptoms of hemolysis | 0
decrease in hemoglobin level | 0
acute renal failure | 0
two sessions of urgent-start hemodialysis | 0
received PRBC | 0
hemolysis attributed to mechanical factors | 0
weak | -720
lethargic | -720
admitted to the hospital | -720
exacerbation of symptoms | -720
hemoglobin level of 6.3 | 0
hematocrit of 19.7 | 0
RBC count of 2.27 | 0
WBC count of 3700 | 0
PLT count of 235000 | 0
MCHC of 32 | 0
MCV of 86.8 | 0
MCH of 27.8 | 0
PT of 15.8 | 0
PTT of 54.4 | 0
INR of 1.2 | 0
Na level of 140 | 0
K level of 4 | 0
BUN of 86 | 0
Cr of 1.3 | 0
uric acid of 9.1 | 0
LDH of 3418 | 0
AST of 64 | 0
ALT of 46 | 0
Alkaline phosphatase of 230 | 0
total bilirubin of 9.6 | 0
direct bilirubin of 2.4 | 0
indirect bilirubin of 7.5 | 0
candidate for blood transfusion | 0
transfusion of first unit of blood initiated | 0
developed fever | 0
developed headache | 0
developed chills | 0
developed back pain | 0
developed urine discoloration | 0
blood transfusion stopped | 0
therapeutic measures taken | 0
blood culture | 0
blood smear | 0
antibody screening test | 0
Coombs test | 0
Coombs Wright test | 0
positive anti-E | 0
positive anti-c | 0
positive anti-Kell | 0
transfused with 3 units of PRBC | 0
ABO compatible | 0
Rh (D) compatible | 0
c-negative | 0
E-negative | 0
Kell-negative | 0
leuko-reduced RBC | 0
Hb raised from 6.3 to 10.5 | 0
transfused 3 more units of PRBC | 0
acceptable Hb level | 0
surgical TV repair | 0
AVR | 0
MVR | 0
transferred to ICU | 0
extubated | 48
no evidence of hemolysis | 48
acceptable Hb level postoperatively | 48
developed sepsis | 504
expired | 504
