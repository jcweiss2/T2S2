32 years old | 0
male | 0
admitted to the hospital | 0
shortness of breath | 0
syncope | 0
seizure | 0
chest pain | 0
flu-like symptoms | -72
intellectual disability | 0
developmental delay | 0
sedentary lifestyle | 0
hypertension | 0
tachycardia | 0
hypotension | 0
hypoxia | 0
oxygen saturation 92% | 0
clear chest auscultation | 0
normal heart sounds | 0
T wave inversions | 0
right ventricular strain | 0
dilated RV | 0
mobile thrombus in right atrium | 0
mobile thrombus in RV | 0
thrombus in transit through PFO | 0
elevated urea | 0
elevated creatinine | 0
high haemoglobin | 0
high haematocrit | 0
dehydration | 0
elevated lactate | 0
elevated D-Dimer | 0
elevated troponin | 0
resuscitation | 0
emergency pulmonary embolectomy | 0
transfer to theatre | 0
prebypass transoesophageal echocardiography | 0
extensive clot in RA | 0
extensive clot in RV | 0
extensive clot in LA | 0
D-shaped septum | 0
severe tricuspid regurgitation | 0
epinephrine infusion | 0
difficulty separating from cardiopulmonary bypass | 0
central ECMO | 0
weaning off CPB | 0
moved to ICU | 0
critical state | 0
full ECMO support | 0
early renal support | 0
continuous venovenous haemodiafiltration | 0
intravenous sildenafil | 0
pulmonary vasodilation | 0
weaning off ECMO | 144
sepsis | 192
acute kidney injury | 192
critical illness neuropathy | 192
aggressive supportive care | 192
respiratory function stabilization | 192
percutaneous tracheostomy | 480
weaning from ventilator | 672
IV heparin | 0
warfarin | 144
oral tadalafil | 144
haematemesis | 720
endoscopy | 720
old traumatic ulcer | 720
clipping of ulcer | 720
tracheostomy tube removal | 888
discharged home | 1032
follow-up outpatient echo | 1008
normalization of RV function | 1008
full recovery | 1008
antinuclear antibodies negative | 0
factor V Leiden mutation negative | 0
anticardiolipin negative | 0
double-stranded DNA antibodies negative | 0
beta-2 glycoprotein-1 antibodies negative | 0
no evidence of Bechet’s disease | 0
no evidence of underlying malignancy | 0
chest CT scan | 0
cytology from bronchoscopy | 0