66 years old | 0
male | 0
diabetes mellitus type 2 | 0
hypertension | 0
dyslipidemia | 0
dry cough | -168
mild shortness of breath | -168
fever | -168
chest X-ray unremarkable | -168
discharged home | -168
RT-PCR positive for SARS-CoV-2 | -168
returned due to worsening shortness of breath | -168
transferred to institution | -168
blood pressure 128/77 mm Hg | 0
heart rate 84 beats/minute | 0
respiratory rate 32 beats/minute | 0
temperature 36.2 °C | 0
oxygen saturation 98% on 6 liters of oxygen | 0
admitted to intensive care unit | 0
treated with hydroxychloroquine | 0
treated with azithromycin | 0
treated with IV ceftriaxone | 0
respiratory distress | 96
severe hypoxia with oxygen saturation of 40% | 96
hemodynamically unstable (blood pressure 50/31 mm Hg) | 96
emergently intubated | 96
resuscitated with 2 liters of IV fluid boluses | 96
required norepinephrine | 96
required vasopressin | 96
required epinephrine infusion | 96
mean arterial pressure above 65 mm Hg | 96
point-of-care cardiac ultrasonography showed severely reduced LVEF | 96
started on dobutamine | 96
arterial blood gas pH 7.17 | 96
arterial blood gas PaCO2 48 | 96
arterial blood gas PaO2 69 | 96
arterial blood gas bicarbonate 19 mmol/L | 96
PaO2/FiO2 ratio of 69 | 96
chest X-ray interval worsening | 96
ECG sinus tachycardia | 96
ECG low voltage complexes | 96
ECG nonspecific T-wave abnormalities | 96
troponin T 0.39 ng/mL | 96
NT-proBNP 798 pg/mL | 96
transthoracic echocardiography severe LV dysfunction | 120
LVEF 32% | 120
global LV hypokinesia | 120
ferritin 100586 ng/mL | 120
lactate dehydrogenase >25000 U/L | 120
D-dimer 6.99 µg/mL | 120
CRP 278.4 mg/L | 120
weaned off norepinephrine | 96
weaned off vasopressin | 96
weaned off epinephrine infusion | 96
supportive treatment mechanical ventilation | 96
supportive treatment antibiotics (IV vancomycin and cefepime) | 96
supportive treatment IV diuretics | 96
convalescent plasma on day 5 | 120
convalescent plasma on day 6 | 144
convalescent plasma on day 12 | 288
cardiogenic shock improved | 192
dobutamine deescalating need | 192
dobutamine discontinued on day 8 | 192
troponin T 0.05 ng/mL | 192
NT-proBNP 26 pg/mL | 192
ferritin 4320 ng/mL | 192
CRP 69.7 mg/L | 192
D-dimer 2.38 µg/mL | 192
LD 427 U/L | 192
repeat transthoracic echocardiography LVEF 60-65% | 240
normal LV systolic function | 240
no wall motion abnormalities | 240
extubated on day 15 | 360
repeat COVID-19 RT-PCR negative | 456
discharged home | 456
