56 years old | 0
male | 0
Malay | 0
admitted to the hospital | 0
abdominal distension | -120
diagnosed with hepatocellular carcinoma | -120
chronic hepatitis B | -120
referred to the institute | -120
dynamic CT scan of the liver | 0
hypervascular lesions at segments IVa, VII and VIII | 0
cirrhosis | 0
splenomegaly | 0
esophageal varices | 0
no ascites | 0
local treatment of the multicentric HCC using RFA | 0
pre-procedural assessment | 0
small ventricular septal defect | 0
left to right shunting | 0
normal chamber sizes | 0
normal left ventricular ejection fraction | 0
Child Class A compensated liver disease | 0
serum albumin 32 g/L | 0
serum bilirubin 21 µmol/L | 0
alanine aminotransferase (ALT) 45 IU/L | 0
aspartate aminotransferase (AST) 54 IU/L | 0
platelet count 61 × 10^9/L | 0
International Normalised Ratio 1.2 | 0
alpha fetoprotein (AFP) 23.8 ng/mL | 0
RFA procedure | 0
general anesthesia | 0
fluoroscopic CT guidance | 0
10 cm long expandable 15 G StarBurst XL radiofrequency (RF) needle | 0
RF current generator | 0
four grounding pads | 0
pulse-oximetry | 0
arterial blood pressure | 0
cardiac activity | 0
CT fluoroscopic guidance | 0
needle tip placement | 0
deployment of thines | 0
ablation of the largest tumour | 0
repositioning of the needle | 0
ablation of the medial and lateral margins | 0
coagulation necrosis | 0
no evidence of any pericardial fluid | 0
difficulty in retracting the thines | 0
haemorrhagic cardiac tamponade | 1
expanding pericardial effusion | 1
pericardiocentesis | 1
haemorrhagic fluid | 1
emergency sternostomy | 2
evacuation of blood from the pericardium | 2
puncture wound at the anterior cardiac vein | 2
inflammatory changes in the adjacent diaphragm | 2
no evidence of any ablation change in the pericardium | 2
repair of the anterior cardiac vein | 2
haemostasis | 2
stable post-surgery | 2
deterioration of condition | 48
liver failure | 48
upper gastrointestinal bleeding | 48
pneumonia | 48
sepsis | 48
expiration | 456
RFA complication | 0
haemorrhagic cardiac tamponade | 1
rare complication | 0
pre-procedural assessment | 0
prevention of complications | 0
early detection | 0
proper management | 0
thermal protection technique | 0
real-time imaging guidance | 0
prevention of charring and tissue adhesion | 0
removal of the RF needle | 0
cleaning and redeployment of the RF needle | 0