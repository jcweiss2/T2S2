There is no time information in the free-form response.