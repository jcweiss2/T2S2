36 years old | 0
female | 0
cerebral palsy | 0
severe kyphoscoliosis | 0
admitted to respiratory intensive care unit | 0
severe respiratory failure | 0
pneumonia | 0
orotracheal intubation | 24
invasive mechanical ventilation | 24
tracheotomy | 168
persistent type II respiratory failure | 168
peristomal skin diastase | 672
tracheocutaneous fistula | 672
excessive cuff pressure | 672
surgical repair | 696
tracheotomy with suturing of the distal stump | 696
surgical treatment | 696
mechanical ventilation through a tracheal cannula | 696
reduced length of the residual trachea | 696
cuff securing system | 696
selective intubation of the main bronchi | 696
inflating the cuffs at both main stem bronchi inlets | 696
Y-shaped bridge | 696
ventilator connection | 696
adequate minute volume | 696
blood gas levels | 696
no significant leaks | 696
ventilatory parameters remained stable | 696
bronchoscopic examination | 700
no evidence of alterations on both main bronchi | 700
died | 736
sepsis | 736