12 years old | 0
neutered female | 0
American cocker spaniel | 0
9.9 kg | 0
BCS 3/5 | 0
admitted to the hospital | 0
dyspnea | -48
anorexia | -48
gallbladder mucocele | -192
pancreatitis | -192
extrahepatic bile duct obstruction | -192
surgically removed | -96
discharged | -96
lethargic | 0
tachypnea | 0
respiratory distress | 0
heart rate 128 bpm | 0
heart murmur not auscultated | 0
SpO2 not measurable | 0
systolic blood pressure 162 mmHg | 0
diastolic blood pressure 69 mmHg | 0
leukocytosis | 0
thrombocytopenia | 0
normal serum biochemical profile | 0
prothrombin time 8.0 sec | 0
activated partial thromboplastin time 21.1 sec | 0
fibrinogen 344 mg/dl | 0
cardiac enlargement | 0
enlargement of the main pulmonary artery | 0
interstitial and alveolar lung patterns | 0
severe RV dilation | 0
right atrial dilation | 0
main PA dilation | 0
myocardial hypokinesis of the RV free wall | 0
interventricular septal flattening | 0
paradoxical septal motion | 0
mild tricuspid regurgitation | 0
high velocity of TR | 0
estimated RA pressure 10 mmHg | 0
estimated systolic PA pressure 93.4 mmHg | 0
asymmetrical PA flow profile | 0
mid-systolic notching | 0
PA acceleration time 35 msec | 0
PA ejection time 204 msec | 0
acceleration time/ejection time ratio 0.17 | 0
impaired relaxation pattern | 0
peak systolic tricuspid annular velocity 10.5 cm/sec | 0
tricuspid annulus plane systolic excursion 7.9 mm | 0
fractional area change 24.7% | 0
Tei index 0.62 | 0
RV free wall longitudinal strain -7.3% | 0
septal longitudinal strain -6.0% | 0
RV-SD 83.4 msec | 0
CT angiography | 0
filling defect in left and right main PA | 0
filling defect in left and right brachiocephalic veins | 0
filling defect in right external jugular vein | 0
atelectasis in the middle lobe | 0
ground-grass opacity in the lung lobes | 0
diagnosed as acute PTE | 0
oxygen therapy initiated | 0
low molecular heparin administered | 0
cefazolin sodium hydrate administered | 0
aspirin administered | 0
clopidogrel sulfate administered | 0
respiratory status improved | 216
breathing normally in room air | 216
echocardiography on day 9 | 216
reduction in the size of the right heart | 216
improvement in interventricular septal flattening | 216
decrease in the velocity of TR | 216
improvement in RV free wall hypokinesis | 216
improvement in RV dyssynchrony | 216
CT angiography on day 9 | 216
filling defects in the PA and brachiocephalic veins unchanged | 216
abnormal findings in lung field disappeared | 216
discharged from hospital | 240
elevated plasma D-dimer | 0
elevated fibrin degradation product | 0