67 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
body weight 50 kg | 0 | 0 | Factual
height 158 cm | 0 | 0 | Factual
backache | -1 | 0 | Factual
calculi in both kidneys | -1 | 0 | Factual
ureteral calculi | -1 | 0 | Factual
admitted to hospital | 0 | 0 | Factual
HLL | 0 | 0 | Factual
double J catheterization | 0 | 0 | Factual
purulent urine | 0 | 0 | Factual
fever | 0.5 | 48 | Factual
chill | 0.5 | 48 | Factual
low blood pressure | 0.5 | 48 | Factual
imipenem and Cilastatin sodium | 0.5 | 48 | Factual
fluid resuscitation | 0.5 | 48 | Factual
Norepinephrine | 0.5 | 48 | Factual
Hydrocortisone sodium succinate | 0.5 | 48 | Factual
anuria | 48 | 48 | Factual
ARDS | 48 | 48 | Factual
invasive ventilatory support | 48 | 240 | Factual
CRRT | 48 | 240 | Factual
transferred to ICU | 48 | 48 | Factual
sedated state | 48 | 48 | Factual
blood pressure 80/62 mmHg | 48 | 48 | Factual
heart rate 139 beats/min | 48 | 48 | Factual
transcutaneous oxygen saturation 80% | 48 | 48 | Factual
cold, clammy extremities | 48 | 48 | Factual
loud bubbling sound in the lung | 48 | 48 | Factual
arterial blood gas analysis | 48 | 48 | Factual
oxygen partial pressure 50 mmHg | 48 | 48 | Factual
lactic acid 10.6 mmol/L | 48 | 48 | Factual
bicarbonate 10.8 mmol/L | 48 | 48 | Factual
central venous pressure 20 cmH2O | 48 | 48 | Factual
B lines in lung ultrasonography | 48 | 48 | Factual
diffuse dysfunction in left ventricle | 48 | 48 | Factual
LVEF 20.3% | 48 | 48 | Factual
normal function in right ventricle | 48 | 48 | Factual
sinus tachycardia | 48 | 48 | Factual
broad ST depression | 48 | 48 | Factual
elevated troponin I | 48 | 48 | Factual
elevated amino-terminal brain natriuretic peptide precursor | 48 | 48 | Factual
creatinine 356 μmol/L | 48 | 48 | Factual
anuria | 48 | 240 | Factual
VA-ECMO | 48 | 144 | Factual
CRRT | 48 | 240 | Factual
imipenem and Cilastatin sodium | 48 | 240 | Factual
Vancomycin | 48 | 240 | Factual
Norepinephrine stopped | 78 | 78 | Factual
Epinephrine stopped | 78 | 78 | Factual
lactic acid level declined | 90 | 90 | Factual
vasoactive drugs stopped | 138 | 138 | Factual
arterial blood lactate level normal | 144 | 144 | Factual
extended-spectrum β-lactamase-positive Escherichia coli | 48 | 48 | Factual
inflammatory indices diminished | 240 | 240 | Factual
anti-infection regimen continued | 240 | 240 | Factual
minimum serum trough concentration of Vancomycin | 240 | 240 | Factual
LVEF 35% | 120 | 120 | Factual
black and necrotic skin | 120 | 120 | Factual
weaned from ECMO | 144 | 144 | Factual
renal function improved | 144 | 144 | Factual
CRRT discontinued | 144 | 144 | Factual
urine volume increased | 144 | 240 | Factual
vascular ultrasonography | 240 | 240 | Factual
computed tomography angiography | 240 | 240 | Factual
vascular surgery consultation | 240 | 240 | Factual
necrotic tissues amputated | 336 | 336 | Factual
respiratory function supported | 48 | 240 | Factual
spontaneous breathing | 120 | 120 | Factual
trachea opened | 240 | 240 | Factual
anti-infective therapy changed | 240 | 240 | Factual
weaned from ventilator | 480 | 480 | Factual
tracheotomy tube sealed | 600 | 600 | Factual
discharged | 768 | 768 | Factual
intermittent hemodialysis | 768 | 768 | Factual
self-care | 1296 | 1296 | Factual
intermittent hemodialysis continued | 1296 | 1296 | Factual