4 years old | 0
male | 0
Saudi | 0
admitted to the hospital | 0
thick platelike hyperkeratotic scales | -672
ectropion | -672
eclabium | -672
harlequin ichthyosis | -672
severe anemia | -672
thrombocytopenia | -672
sepsis | -672
skin care | -672
desquamated | -56
well-demarcated symmetric erythematous thick hyperkeratotic plaques | -56
fixed flexion deformity of the elbows | -56
fixed flexion deformity of the hands | -56
fixed flexion deformity of the feet | -56
mitten hand deformity | -56
sharply demarcated erythematous scaly plaque | -56
whole-exome sequencing | -56
whole-genome sequencing | -56
homozygous missense variant in KDSR | -56
novel homozygous variant | -56
skeletal surveys | -56
bone marrow biopsy | -56
congenital megakaryocytic aplasia | -56
skin biopsy | -56
nonspecific hyperkeratosis | -56
acanthosis | -56
papillary dermis fibrosis | -56
discharged | 56
sepsis | 120
epistaxis | 120
mild subdural hematoma | 120
platelet transfusions | 120
intravenous immunoglobulin | 120
packed red blood cells | 120
acitretin | 120
isotretinoin | 240
good control of skin condition | 240
flareups during febrile episodes | 240 
death of sister | -8760
cesarean section | -672 
consanguineous parents | 0 
elective birth | -672 
transport to tertiary center | -656 
admitted to neonatal intensive care unit | -672 
multiple transfusions | -672 
intravenous antibiotics | -672 
recurrent sepsis | -672 
thick scales | -672 
gradual desquamation | -56 
erythematous scaly plaque | -56 
upper half of face | -56 
erythrokeratodermas | 0 
autosomal dominant | 0 
autosomal recessive | 0 
genetic skin disorders | 0 
well-demarcated symmetric thick plaques | 0 
variable clinical pictures | 0 
focal red hyperkeratotic plaques | 0 
palmoplantar scaling | 0 
collodion membrane | 0 
thrombocytopenia | 0 
anemia | 0 
platelet counts | 120 
hemoglobin levels | 120 
retinoic acid derivatives | 240 
sphingosine acylation | 240 
sphingomyelinase | 240 
de novo pathway | 240 
KDSR mutations | 0 
broad spectrum of clinical manifestations | 0 
HI-like features | 0 
localized keratodermas | 0 
severe self-resolving hematological manifestations | 0 
persistent hematological manifestations | 0 
novel variant | 0 
long-term sequelae | 0 
prognosis | 0 
survival | 0 
close monitoring | 0 
differential diagnosis | 0 
pathogenesis of non-ABCA12 HI | 0 
ABCA12 gene mutations | 0 
harlequin ichthyosis | 0 
harlequin phenotype | 0 
erythroderma | 0 
small scales | 0 
neonates | 0 
rare genetic skin disorders | 0 
Progressive symmetrical erythrokeratoderma | 0 
PSEK | 0 
Gottron syndrome | 0 
fixed symmetric well-demarcated hyperkeratotic plaques | 0 
peripheral erythema | 0 
extensor surfaces | 0 
face | 0 
trunk | 0 
homozygous variant | 0 
KDSR gene | 0 
3-ketodihydrosphingosine reductase | 0 
whole-genome sequencing | 0 
NM_002035.4:c.434A>G | 0 
p. Asn145Ser | 0 
gnomAD | 0 
local database | 0 
in silico tools | 0 
CADD | 0 
DANN | 0 
PolyPhen | 0 
SIFT | 0 
GERP | 0 
pathogenic | 0 
clinical picture | 0 
thick plates | 0 
erythroderma | 0 
fine scales | 0 
spontaneous resolution | 0 
persistent severe thrombocytopenia | 0 
hepatic hemangioendothelioma | 0 
de novo synthesis pathway | 0 
sphingolipids | 0 
megakaryopoiesis | 0 
cytoplasmic organization | 0 
proplatelet formation | 0 
skin integrity | 0 
cutaneous proliferation | 0 
differentiation | 0 
perturbation | 0 
sphingosine acylation | 0 
sphingomyelinase | 0 
independent pathways | 0 
retinoic acid derivatives | 0 
near-complete resolution | 0 
up-regulation | 0 
sphingomyelinase | 0 
independent of the de novo pathway | 0 
broad spectrum of clinical manifestations | 0 
HI-like features | 0 
localized keratodermas | 0 
severe self-resolving hematological manifestations | 0 
persistent hematological manifestations | 0 
novel variant | 0 
long-term sequelae | 0 
prognosis | 0 
survival | 0 
close monitoring | 0 
differential diagnosis | 0 
pathogenesis of non-ABCA12 HI | 0 
ABCA12 gene mutations | 0 
harlequin ichthyosis | 0 
harlequin phenotype | 0 
erythroderma | 0 
small scales | 0 
neonates | 0 
rare genetic skin disorders | 0 
Progressive symmetrical erythrokeratoderma | 0 
PSEK | 0 
Gottron syndrome | 0 
fixed symmetric well-demarcated hyperkeratotic plaques | 0 
peripheral erythema | 0 
extensor surfaces | 0 
face | 0 
trunk | 0 
homozygous variant | 0 
KDSR gene | 0 
3-ketodihydrosphingosine reductase | 0 
whole-genome sequencing | 0 
NM_002035.4:c.434A>G | 0 
p. Asn145Ser | 0 
gnomAD | 0 
local database | 0 
in silico tools | 0 
CADD | 0 
DANN | 0 
PolyPhen | 0 
SIFT | 0 
GERP | 0 
pathogenic | 0 
clinical picture | 0 
thick plates | 0 
erythroderma | 0 
fine scales | 0 
spontaneous resolution | 0 
persistent severe thrombocytopenia | 0 
hepatic hemangioendothelioma | 0 
de novo synthesis pathway | 0 
sphingolipids | 0 
megakaryopoiesis | 0 
cytoplasmic organization | 0 
proplatelet formation | 0 
skin integrity | 0 
cutaneous proliferation | 0 
differentiation | 0 
perturbation | 0 
sphingosine acylation | 0 
sphingomyelinase | 0 
independent pathways | 0 
retinoic acid derivatives | 0 
near-complete resolution | 0 
up-regulation | 0 
sphingomyelinase | 0 
independent of the de novo pathway | 0 
broad spectrum of clinical manifestations | 0 
HI-like features | 0 
localized keratodermas | 0 
severe self-resolving hematological manifestations | 0 
persistent hematological manifestations | 0 
novel variant | 0 
long-term sequelae | 0 
prognosis | 0 
survival | 0 
close monitoring | 0 
differential diagnosis | 0 
pathogenesis of non-ABCA12 HI | 0 
ABCA12 gene mutations | 0 
harlequin ichthyosis | 0 
harlequin phenotype | 0 
erythroderma | 0 
small scales | 0 
neonates | 0 
rare genetic skin disorders | 0 
Progressive symmetrical erythrokeratoderma | 0 
PSEK | 0 
Gottron syndrome | 0 
fixed symmetric well-demarcated hyperkeratotic plaques | 0 
peripheral erythema | 0 
extensor surfaces | 0 
face | 0 
trunk | 0 
homozygous variant | 0 
KDSR gene | 0 
3-ketodihydrosphingosine reductase | 0 
whole-genome sequencing | 0 
NM_002035.4:c.434A>G | 0 
p. Asn145Ser | 0 
gnomAD | 0 
local database | 0 
in silico tools | 0 
CADD | 0 
DANN | 0 
PolyPhen | 0 
SIFT | 0 
GERP | 0 
pathogenic | 0 
clinical picture | 0 
thick plates | 0 
erythroderma | 0 
fine scales | 0 
spontaneous resolution | 0 
persistent severe thrombocytopenia | 0 
hepatic hemangioendothelioma | 0 
de novo synthesis pathway | 0 
sphingolipids | 0 
megakaryopoiesis | 0 
cytoplasmic organization | 0 
proplatelet formation | 0 
skin integrity | 0 
cutaneous proliferation | 0 
differentiation | 0 
perturbation | 0 
sphingosine acylation | 0 
sphingomyelinase | 0 
independent pathways | 0 
retinoic acid derivatives | 0 
near-complete resolution | 0 
up-regulation | 0 
sphingomyelinase | 0 
independent of the de novo pathway | 0 
broad spectrum of clinical manifestations | 0 
HI-like features | 0 
localized keratodermas | 0 
severe self-resolving hematological manifestations | 0 
persistent hematological manifestations | 0 
novel variant | 0 
long-term sequelae | 0 
prognosis | 0 
survival | 0 
close monitoring | 0 
differential diagnosis | 0 
pathogenesis of non-ABCA12 HI | 0 
ABCA12 gene mutations | 0 
harlequin ichthyosis | 0 
harlequin phenotype | 0 
erythroderma | 0 
small scales | 0 
neonates | 0 
rare genetic skin disorders | 0 
Progressive symmetrical erythrokeratoderma | 0 
PSEK | 0 
Gottron syndrome | 0 
fixed symmetric well-demarcated hyperkeratotic plaques | 0 
peripheral erythema | 0 
extensor surfaces | 0 
face | 0 
trunk | 0 
homozygous variant | 0 
KDSR gene | 0 
3-ketodihydrosphingosine reductase | 0 
whole-genome sequencing | 0 
NM_002035.4:c.434A>G | 0 
p. Asn145Ser | 0 
gnomAD | 0 
local database | 0 
in silico tools | 0 
CADD | 0 
DANN | 0 
PolyPhen | 0 
SIFT | 0 
GERP | 0 
pathogenic | 0 
clinical picture | 0 
thick plates | 0 
erythroderma | 0 
fine scales | 0 
spontaneous resolution | 0 
persistent severe thrombocytopenia | 0 
hepatic hemangioendothelioma | 0 
de novo synthesis pathway | 0 
sphingolipids | 0 
megakaryopoiesis | 0 
cytoplasmic organization | 0 
proplatelet formation | 0 
skin integrity | 0 
cutaneous proliferation | 0 
differentiation | 0 
perturbation | 0 
sphingosine acylation | 0 
sphingomyelinase | 0 
independent pathways | 0 
retinoic acid derivatives | 0 
near-complete resolution | 0 
up-regulation | 0 
sphingomyelinase | 0 
independent of the de novo pathway | 0 
broad spectrum of clinical manifestations | 0 
HI-like features | 0 
localized keratodermas | 0 
severe self-resolving hematological manifestations | 0 
persistent hematological manifestations | 0 
novel variant | 0 
long-term sequelae | 0 
prognosis | 0 
survival | 0 
close monitoring | 0 
differential diagnosis | 0 
pathogenesis of non-ABCA12 HI | 0 
ABCA12 gene mutations | 0 
harlequin ichthyosis | 0 
harlequin phenotype | 0 
erythroderma | 0 
small scales | 0 
neonates | 0 
rare genetic skin disorders | 0 
Progressive symmetrical erythrokeratoderma | 0 
PSEK | 0 
Gottron syndrome | 0 
fixed symmetric well-demarcated hyperkeratotic plaques | 0 
peripheral erythema | 0 
extensor surfaces | 0 
face | 0 
trunk | 0 
homozygous variant | 0 
KDSR gene | 0 
3-ketodihydrosphingosine reductase | 0 
whole-genome sequencing | 0 
NM_002035.4:c.434A>G | 0 
p. Asn145Ser | 0 
gnomAD | 0 
local database | 0 
in silico tools | 0 
CADD | 0 
DANN | 0 
PolyPhen | 0 
SIFT | 0 
GERP | 0 
pathogenic | 0 
clinical picture | 0 
thick plates | 0 
erythroderma | 0 
fine scales | 0 
spontaneous resolution | 0 
persistent severe thrombocytopenia | 0 
hepatic hemangioendothelioma | 0 
de novo synthesis pathway | 0 
sphingolipids | 0 
megakaryopoiesis | 0 
cytoplasmic organization | 0 
proplatelet formation | 0 
skin integrity | 0 
cutaneous proliferation | 0 
differentiation | 0 
perturbation | 0 
sphingosine acylation | 0 
sphingomyelinase | 0 
independent pathways | 0 
retinoic acid derivatives | 0 
near-complete resolution | 0 
up-regulation | 0 
sphingomyelinase | 0 
independent of the de novo pathway | 0 
broad spectrum of clinical manifestations | 0 
HI-like features | 0 
localized keratodermas | 0 
severe self-resolving hematological manifestations | 0 
persistent hematological manifestations | 0 
novel variant | 0 
long-term sequelae | 0 
prognosis | 0 
survival | 0 
close monitoring | 0 
differential diagnosis | 0 
pathogenesis of non-ABCA12 HI | 0 
ABCA12 gene mutations | 0 
harlequin ichthyosis | 0 
harlequin phenotype | 0 
erythroderma | 0 
small scales | 0 
neonates | 0 
rare genetic skin disorders | 0 
Progressive symmetrical erythrokeratoderma | 0 
PSEK | 0 
Gottron syndrome | 0 
fixed symmetric well-demarcated hyperkeratotic plaques | 0 
peripheral erythema | 0 
extensor surfaces | 0 
face | 0 
trunk | 0 
homozygous variant | 0 
KDSR gene | 0 
3-ketodihydrosphingosine reductase | 0 
whole-genome sequencing | 0 
NM_002035.4:c.434A>G | 0 
p. Asn145Ser | 0 
gnomAD | 0 
local database | 0 
in silico tools | 0 
CADD | 0 
DANN | 0 
PolyPhen | 0 
SIFT | 0 
GERP | 0 
pathogenic | 0 
clinical picture | 0 
thick plates | 0 
erythroderma | 0 
fine scales | 0 
spontaneous resolution | 0 
persistent severe thrombocytopenia | 0 
hepatic hemangioendothelioma | 0 
de novo synthesis pathway | 0 
sphingolipids | 0 
megakaryopoiesis | 0 
cytoplasmic organization | 0 
proplatelet formation | 0 
skin integrity | 0 
cutaneous proliferation | 0 
differentiation | 0 
perturbation | 0 
sphingosine acylation | 0 
sphingomyelinase | 0 
independent pathways | 0 
retinoic acid derivatives | 0 
near-complete resolution | 0 
up-regulation | 0 
sphingomyelinase | 0 
independent of the de novo pathway | 0 
broad spectrum of clinical manifestations | 0 
HI-like features | 0 
localized keratodermas | 0 
severe self-resolving hematological manifestations | 0 
persistent hematological manifestations | 0 
novel variant | 0 
long-term sequelae | 0 
prognosis | 0 
survival | 0 
close monitoring | 0 
differential diagnosis | 0 
pathogenesis of non-ABCA12 HI | 0 
ABCA12 gene mutations | 0 
harlequin ichthyosis | 0 
harlequin phenotype | 0 
erythroderma | 0 
small scales | 0 
neonates | 0 
rare genetic skin disorders | 0 
Progressive symmetrical erythrokeratoderma | 0 
PSEK | 0 
Gottron syndrome | 0 
fixed symmetric well-demarcated hyperkeratotic plaques | 0 
peripheral erythema | 0 
extensor surfaces | 0 
face | 0 
trunk | 0 
homozygous variant | 0 
KDSR gene | 0 
3-ketodihydrosphingosine reductase | 0 
whole-genome sequencing | 0 
NM_002035.4:c.434A>G | 0 
p. Asn145Ser | 0 
gnomAD | 0 
local database | 0 
in silico tools | 0 
CADD | 0 
DANN | 0 
PolyPhen | 0 
SIFT | 0 
GERP | 0 
pathogenic | 0 
clinical picture | 0 
thick plates | 0 
erythroderma | 0 
fine scales | 0 
spontaneous resolution | 0 
persistent severe thrombocytopenia | 0 
hepatic hemangioendothelioma | 0 
de novo synthesis pathway | 0 
sphingolipids | 0 
megakaryopoiesis | 0 
cytoplasmic organization | 0 
proplatelet formation | 0 
skin integrity | 0 
cutaneous proliferation | 0 
differentiation | 0 
perturbation | 0 
sphingosine acylation | 0 
sphingomyelinase | 0 
independent pathways | 0 
retinoic acid derivatives | 0 
near-complete resolution | 0 
up-regulation | 0 
sphingomyelinase | 0 
independent of the de novo pathway | 0 
broad spectrum of clinical manifestations | 0 
HI-like features | 0 
localized keratodermas | 0 
severe self-resolving hematological manifestations | 0 
persistent hematological manifestations | 0 
novel variant | 0 
long-term sequelae | 0 
prognosis | 0 
survival | 0 
close monitoring | 0 
differential diagnosis | 0 
pathogenesis of non-ABCA12 HI | 0 
ABCA12 gene mutations | 0 
harlequin ichthyosis | 0 
harlequin phenotype | 0 
erythroderma | 0 
small scales | 0 
neonates | 0 
rare genetic skin disorders | 0 
Progressive symmetrical erythrokeratoderma | 0 
PSEK | 0 
Gottron syndrome | 0 
fixed symmetric well-demarcated hyperkeratotic plaques | 0 
peripheral erythema | 0 
extensor surfaces | 0 
face | 0 
trunk | 0 
homozygous variant | 0 
KDSR gene | 0 
3-ketodihydrosphingosine reductase | 0 
whole-genome sequencing | 0 
NM_002035.4:c.434A>G | 0 
p. Asn145Ser | 0 
gnomAD | 0 
local database | 0 
in silico tools | 0 
CADD | 0 
DANN | 0 
PolyPhen | 0 
SIFT | 0 
GERP | 0 
pathogenic | 0 
clinical picture | 0 
thick plates | 0 
erythroderma | 0 
fine scales | 0 
spontaneous resolution | 0 
persistent severe thrombocytopenia | 0 
hepatic hemangioendothelioma | 0 
de novo synthesis pathway | 0 
sphingolipids | 0 
megakaryopoiesis | 0 
cytoplasmic organization | 0 
proplatelet formation | 0 
skin integrity | 0 
cutaneous proliferation | 0 
differentiation | 0 
perturbation | 0 
sphingosine acylation | 0 
sphingomyelinase | 0 
independent pathways | 0 
retinoic acid derivatives | 0 
near-complete resolution | 0 
up-regulation | 0 
sphingomyelinase | 0 
independent of the de novo pathway | 0 
broad spectrum of clinical manifestations | 0 
HI-like features | 0 
localized keratodermas | 0 
severe self-resolving hematological manifestations | 0 
persistent hematological manifestations | 0 
novel variant | 0 
long-term sequelae | 0 
prognosis | 0 
survival | 0 
close monitoring | 0 
differential diagnosis | 0 
pathogenesis of non-ABCA12 HI | 0 
ABCA12 gene mutations | 0 
harlequin ichthyosis | 0 
harlequin phenotype | 0 
erythroderma | 0 
small scales | 0 
neonates | 0 
rare genetic skin disorders | 0 
Progressive symmetrical erythrokeratoderma | 0 
PSEK | 0 
Gottron syndrome | 0 
fixed symmetric well-demarcated hyperkeratotic plaques | 0 
peripheral erythema | 0 
extensor surfaces | 0 
face | 0 
trunk | 0 
homozygous variant | 0 
KDSR gene | 0 
3-ketodihydrosphingosine reductase | 0 
whole-genome sequencing | 0 
NM_002035.4:c.434A>G | 0 
p. Asn145Ser | 0 
gnomAD | 0 
local database | 0 
in silico tools | 0 
CADD | 0 
DANN | 0 
PolyPhen | 0 
SIFT | 0 
GERP | 0 
pathogenic | 0 
clinical picture | 0 
thick plates | 0 
erythroderma | 0 
fine scales | 0 
spontaneous resolution | 0 
persistent severe thrombocytopenia | 0 
hepatic hemangioendothelioma | 0 
de novo synthesis pathway | 0 
sphingolipids | 0 
megakaryopoiesis | 0 
cytoplasmic organization | 0 
proplatelet formation | 0 
skin integrity | 0 
cutaneous proliferation | 0 
differentiation | 0 
perturbation | 0 
sphingosine acylation | 0 
sphingomyelinase | 0 
independent pathways | 0 
retinoic acid derivatives | 0 
near-complete resolution | 0 
up-regulation | 0 
sphingomyelinase | 0 
independent of the de novo pathway | 0 
broad spectrum of clinical manifestations | 0 
HI-like features | 0 
localized keratodermas | 0 
severe self-resolving hematological manifestations | 0 
persistent hematological manifestations | 0 
novel variant | 0 
long-term sequelae | 0 
prognosis | 0 
survival | 0 
close monitoring | 0 
differential diagnosis | 0 
pathogenesis of non-ABCA12 HI | 0 
ABCA12 gene mutations | 0 
harlequin ichthyosis | 0 
harlequin phenotype | 0 
erythroderma | 0 
small scales | 0 
neonates | 0 
rare genetic skin disorders | 0 
Progressive symmetrical erythrokeratoderma | 0 
PSEK | 0 
Gottron syndrome | 0 
fixed symmetric well-demarcated hyperkeratotic plaques | 0 
peripheral erythema | 0 
extensor surfaces | 0 
face | 0 
trunk | 0 
homozygous variant | 0 
KDSR gene | 0 
3-ketodihydrosphingosine reductase | 0 
whole-genome sequencing | 0 
NM_002035.4:c.434A>G | 0 
p. Asn145Ser | 0 
gnomAD | 0 
local database | 0 
in silico tools | 0 
CADD | 0 
DANN | 0 
PolyPhen | 0 
SIFT | 0 
GERP | 0 
pathogenic | 0 
clinical picture | 0 
thick plates | 0 
erythroderma | 0 
fine scales | 0 
spontaneous resolution | 0 
persistent severe thrombocytopenia | 0 
hepatic hemangioendothelioma | 0 
de novo synthesis pathway | 0 
sphingolipids | 0 
megakaryopoiesis | 0 
cytoplasmic organization | 0 
proplatelet formation | 0 
skin integrity | 0 
cutaneous proliferation | 0 
differentiation | 0 
perturbation | 0 
sphingosine acylation | 0 
sphingomyelinase | 0 
independent pathways | 0 
retinoic acid derivatives | 0 
near-complete resolution | 0 
up-regulation | 0 
sphingomyelinase | 0 
independent of the de novo pathway | 0 
broad spectrum of clinical manifestations | 0 
HI-like features | 0 
localized keratodermas | 0 
severe self-resolving hematological manifestations | 0 
persistent hematological manifestations | 0 
novel variant | 0 
long-term sequelae | 0 
prognosis | 0 
survival | 0 
close monitoring | 0 
differential diagnosis | 0 
pathogenesis of non-ABCA12 HI | 0 
ABCA12 gene mutations | 0 
harlequin ichthyosis | 0 
harlequin phenotype | 0 
erythroderma | 0 
small scales | 0 
neonates | 0 
rare genetic skin disorders | 0 
Progressive symmetrical erythrokeratoderma | 0 
PSEK | 0 
Gottron syndrome | 0 
fixed symmetric well-demarcated hyperkeratotic plaques | 0 
peripheral erythema | 0 
extensor surfaces | 0 
face | 0 
trunk | 0 
homozygous variant | 0 
KDSR gene | 0 
3-ketodihydrosphingosine reductase | 0 
whole-genome sequencing | 0 
NM_002035.4:c.434A>G | 0 
p. Asn145Ser | 0 
gnomAD | 0 
local database | 0 
in silico tools | 0 
CADD | 0 
DANN | 0 
PolyPhen | 0 
SIFT | 0 
GERP | 0 
pathogenic | 0 
clinical picture | 0 
thick plates | 0 
erythroderma | 0 
fine scales | 0 
spontaneous resolution | 0 
persistent severe thrombocytopenia | 0 
hepatic hemangioendothelioma | 0 
de novo synthesis pathway | 0 
sphingolipids | 0 
megakaryopoiesis | 0 
cytoplasmic organization | 0 
proplatelet formation | 0 
skin integrity | 0 
cutaneous proliferation | 0 
differentiation | 0 
perturbation | 0 
sphingosine acylation | 0 
sphingomyelinase | 0 
independent pathways | 0 
retinoic acid derivatives | 0 
near-complete resolution | 0 
up-regulation | 0 
sphingomyelinase | 0 
independent of the de novo pathway | 0 
broad spectrum of clinical manifestations | 0 
HI-like features | 0 
localized keratodermas | 0 
severe self-resolving hematological manifestations | 0 
persistent hematological manifestations | 0 
novel variant | 0 
long-term sequelae | 0 
prognosis | 0 
survival | 0 
close monitoring | 0 
differential diagnosis | 0 
pathogenesis of non-ABCA12 HI | 0 
ABCA12 gene mutations | 0 
harlequin ichthyosis | 0 
harlequin phenotype | 0 
erythroderma | 0 
small scales | 0 
neonates | 0 
rare genetic skin disorders | 0 
Progressive symmetrical erythrokeratoderma | 0 
PSEK | 0 
Gottron syndrome | 0 
fixed symmetric well-demarcated hyperkeratotic plaques | 0 
peripheral erythema | 0 
extensor surfaces | 0 
face | 0 
trunk | 0 
homozygous variant | 0 
KDSR gene | 0 
3-ketodihydrosphingosine reductase | 0 
whole-genome sequencing | 0 
NM_002035.4:c.434A>G | 0 
p. Asn145Ser | 0 
gnomAD | 0 
local database | 0 
in silico tools | 0 
CADD | 0 
DANN | 0 
PolyPhen | 0 
SIFT | 0 
GERP | 0 
pathogenic | 0 
clinical picture | 0 
thick plates | 0 
erythroderma | 0 
fine scales | 0 
spontaneous resolution | 0 
persistent severe thrombocytopenia | 0 
hepatic hemangioendothelioma | 0 
de novo synthesis pathway | 0 
sphingolipids | 0 
megakaryopoiesis | 0 
cytoplasmic organization | 0 
proplatelet formation | 0 
skin integrity | 0 
cutaneous proliferation | 0 
differentiation | 0 
perturbation | 0 
sphingosine acylation | 0 
sphingomyelinase | 0 
independent pathways | 0 
retinoic acid derivatives | 0 
near-complete resolution | 0 
up-regulation | 0 
sphingomyelinase | 0 
independent of the de novo pathway | 0 
broad spectrum of clinical manifestations | 0 
HI-like features | 0 
localized keratodermas | 0 
severe self-resolving hematological manifestations | 0 
persistent hematological manifestations | 0 
novel variant | 0 
long-term sequelae | 0 
prognosis | 0 
survival | 0 
close monitoring | 0 
differential diagnosis | 0 
pathogenesis of non-ABCA12 HI | 0 
ABCA12 gene mutations | 0 
harlequin ichthyosis | 0 
harlequin phenotype | 0 
erythroderma | 0 
small scales | 0 
neonates | 0 
rare genetic skin disorders | 0 
Progressive symmetrical erythrokeratoderma | 0 
PSEK | 0 
Gottron syndrome | 0 
fixed symmetric well-demarcated hyperkeratotic plaques | 0 
peripheral erythema | 0 
extensor surfaces | 0 
face | 0 
trunk | 0 
homozygous variant | 0 
KDSR gene | 0 
3-ketodihydrosphingosine reductase | 0 
whole-genome sequencing | 0 
NM_002035.4:c.434A>G | 0 
p. Asn145Ser | 0 
gnomAD | 0 
local database | 0 
in silico tools | 0 
CADD | 0 
DANN | 0 
PolyPhen | 0 
SIFT | 0 
GERP | 0 
pathogenic | 0 
clinical picture | 0 
thick plates | 0 
erythroderma | 0 
fine scales | 0 
spontaneous resolution | 0 
persistent severe thrombocytopenia | 0 
hepatic hemangioendothelioma | 0 
de novo synthesis pathway | 0 
sphingolipids | 0 
megakaryopoiesis | 0 
cytoplasmic organization | 0 
proplatelet formation | 0 
skin integrity | 0 
cutaneous proliferation | 0 
differentiation | 0 
perturbation | 0 
sphingosine acylation | 0 
sphingomyelinase | 0 
independent pathways | 0 
retinoic acid derivatives | 0 
near-complete resolution | 0 
up-regulation | 0 
sphingomyelinase | 0 
independent of the de novo pathway | 0 
broad spectrum of clinical manifestations | 0 
HI-like features | 0 
localized keratodermas | 0 
severe self-resolving hematological manifestations | 0 
persistent hematological manifestations | 0 
novel variant | 0 
long-term sequelae | 0 
prognosis | 0 
survival | 0 
close monitoring | 0 
differential diagnosis | 0 
pathogenesis of non-ABCA12 HI | 0 
ABCA12 gene mutations | 0 
harlequin ichthyosis | 0 
harlequin phenotype | 0 
erythroderma | 0 
small scales | 0 
neonates | 0 
rare genetic skin disorders | 0