83 years old | 0
    male | 0
    admitted to the hospital | 0
    disorientation | 0
    weakness | 0
    went out into the cold | -24
    developed a terrible cough | -24
    treated with GnRH agonist (leuprolide acetate) | -5808
    prostate cancer | -5808
    living independently | -5808
    working as a stonemason | -5808
    began to notice fatigue | -2160
    itching | -2160
    cold intolerance | -2160
    whole-body edema | -2160
    medications included bicalutamide | 0
    silodosin | 0
    antihistamine | -168
    pruritus | -168
    medical history of tuberculosis | 0
    thyroid function not assessed previously | 0
    no abnormal findings indicating hypothyroidism | 0
    sons taking levothyroxine for Hashimoto's disease | 0
    pale appearance | 0
    depressed level of consciousness (GCS 9) | 0
    blood pressure 77/44 mmHg | 0
    pulse 37 beats/min | 0
    axillary body temperature 34.2℃ | 0
    respiratory rate 20 breaths/min | 0
    oxygen saturation 98% | 0
    distant heart sounds | 0
    regular heart rhythm | 0
    decreased breath sounds | 0
    thyroid not palpable | 0
    sparse hair | 0
    thinning of the outer eyebrows | 0
    macroglossia | 0
    hoarse voice | 0
    thickened skin | 0
    marked hyperkeratosis | 0
    profound pitting edema in lower extremities | 0
    increased aspartate transaminase | 0
    increased creatine kinase | 0
    increased brain natriuretic peptide | 0
    no elevations in cardiac enzymes | 0
    sinus bradycardia | 0
    low voltage on ECG | 0
    chest X-ray showed cardiomegaly | 0
    echocardiogram showed normal cardiac structure | 0
    transferred to ICU | 0
    diagnosed with sick sinus syndrome | 0
    started on catecholamines infusion | 0
    pulse rate increased to 50 beats/min | 24
    blood pressure 90/40 mmHg | 24
    persistent impaired consciousness | 24
    hypothermia (34.5℃) | 24
    elevated TSH (76.01 μIU/mL) | 24
    low free T4 (<0.40 ng/dL) | 24
    low free T3 (1.05 pg/mL) | 24
    high anti-thyroid antibodies | 24
    thyroid ultrasonography showed atrophic gland | 24
    diagnosis of myxedema coma | 0
    oral administration of levothyroxine | 0
    oral administration of levotriiodothyronin | 0
    hemodynamics improved | 72
    withdrawal of catecholamine infusion | 72
    consciousness deteriorated to coma | 72
    endotracheal intubation | 72
    shock state (50/30 mmHg) | 72
    continued thyroid hormone replacement | 72
    LT4 via nasogastric tube | 72
    LT3 via nasogastric tube | 72
    additional LT4 via suppository | 72
    elevation in free T4 and T3 levels | 120
    general condition improved | 120
    withdrawal hypothermia | 120
    discontinued catecholamine infusion | 144
    sedative agent given for body motion | 168
    recombinant human thrombomodulin administered | 168
    regained full consciousness | 264
    discharged from ICU | 264
    extubation performed | 360
    relapse of hypercapnia | 360
    placed on NIPPV | 360
    whole-body computed tomography performed | 360
    swelling of the pancreas | 360
    mesenteric edema | 360
    effusion | 360
    fat stranding | 360
    acute pancreatitis | 360
    amylase level 566 IU/L on day 3 | 72
    tube feeding started | 360
    respiratory rehabilitation | 360
    sudden abdominal pain on day 33 | 792
    CT showed increased peripancreatic effusion | 792
    fibrous capsule formation | 792
    elevated WBC (27,200/μL) | 792
    elevated CRP (14.38 mg/dL) | 792
    no elevation of pancreatic enzymes | 792
    possible secondary infection | 792
    broad-spectrum antibiotics administered | 792
    septic shock | 840
    died | 840
    autopsy showed pancreatic necrosis | 840
    retroperitoneal abscesses | 840
    diffuse inflammatory changes in pancreas | 840
    atrophic thyroid with Hashimoto's thyroiditis | 840
    reduction in prostate cancer | 840