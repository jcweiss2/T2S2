59 years old | 0
male | 0
sudden chest pain | -24
collapsed in the ambulance | -24
ventricular fibrillation | -24
cardiopulmonary resuscitation | -24
return of spontaneous circulation | -24
blood pressure 105/78 mm Hg | 0
heart rate 120 beats/min | 0
respiratory rate 20 breaths/min | 0
body temperature 35.8°C | 0
ST-segment elevation myocardial infarction | 0
repeated cardiac arrest | 0
veno-arterial ECMO | 0
percutaneous coronary intervention | 0
thrombectomy | 0
admitted to ICU | 0
sedation with remifentanil | 0
propofol infusion | 0
hemodynamic status improved | 72
oxygenation improved | 72
VA ECMO decannulation | 72
progressive acute kidney injury | 168
continuous renal replacement therapy | 168
severe acute respiratory distress syndrome | 192
hospital-acquired pneumonia | 192
venoCvenous ECMO | 192
clinical improvement of pneumonia | 384
VV ECMO weaned off | 384
sedation retained | 432
vasopressors tapered | 432
increased alanine aminotransferase | 432
increased aspartate aminotransferase | 432
bundle branch block | 480
increased creatinine kinase | 480
increased CK-MB | 480
increased troponin I | 480
aggravated hypotension | 480
increased norepinephrine | 480
increased epinephrine | 480
vasopressin added | 480
acute renal failure | 480
metabolic acidosis | 480
propofol administration | 0
discontinuation of propofol | 504
serum triglyceride level 369 mg/dl | 504
normal cortisol level | 504
normal thyroid function tests | 504
vasopressors requirement decreased | 528
vasopressin tapered | 528
CK level continued to elevate | 528
L-carnitine administration | 552
CK level decline | 648
stabilized with low-dose norepinephrine | 648
discharged from ICU | 1224
transferred to nursing hospital | 2208
lactic acidosis | 480
rhabdomyolysis | 480
arrhythmia | 480
unstable hemodynamics | 480
PRIS diagnosis | 504
no metabolic acidosis | 480
no hyperkalemia | 480
increased lactic acid | 480
elevated CK | 480
elevated myoglobin | 480
hyperlipidemia | 480
ECG changes | 480
masked metabolic acidosis | 480
masked rhabdomyolysis | 480
increased energy demand | 480
decreased energy availability | 480
depletion of ATP | 480
cellular hypoxia | 480
decreased cardiac function | 480
resistance to inotropes | 480
high cumulative propofol dose | 504
high-dose vasopressors | 504
sepsis | 480
neurological injuries | 480
catecholamine use | 480
glucocorticoid use | 480
carbohydrate exhaustion | 480
carnitine deficiency | 480
inborn impairment of fatty acid oxidation | 480
critical illness | 480
ECMO implementation | 480
CRRT application | 480
ventilator synchrony issues | 480
agitation | 480
ventilator dyssynchrony | 480
low-dose propofol infusion | 0
prolonged propofol administration | 504
multimodal sedation regimen | 504
alternative sedatives | 504
PH monitoring | 504
lactate monitoring | 504
triglyceride monitoring | 504
CK monitoring | 504
cardiac marker monitoring | 504
carbohydrate supplementation | 504
lipid minimization | 504
L-carnitine effect uncertain | 552
favorable outcome | 2208
