18 years old | 0
female | 0
admitted to the hospital | 0
increasing abdominal pain | -72
frequency of uterine contractions | -72
intensity of uterine contractions | -72
suprapubic pain | -72
urinary discomfort | -72
vaginal discharge | -72
seen 3 days prior | -72
abnormal vaginal discharge | -72
low abdominal pain | -72
positive fetal fibronectin test | -72
risk of preterm labor | -72
no rupture of membranes | -72
discharged | -72
expectant management | -72
instructed to present to Arnot Ogden Medical Center | -72
prematurity | -72
increase in uterine contractions | -72
past medical history of seizures | -672
past medical history of depression | -672
not currently on medication | 0
remote history of smoking | -6720
respiratory symptoms | -168
shortness of breath | -168
coughing | -168
rhinorrhea | -168
instructed to use over-the-counter medications | -72
symptomatic relief | -72
told symptoms would resolve on own | -72
presumably viral illness | -72
previously living in water-damaged place | -336
utilizing a humidifier | -336
moved out 1 week prior | -168
G1P0 | 0
34 weeks 6 days | 0
routine prenatal care | 0
consistent prenatal care | 0
non-completion of glucose tolerance test | 0
remained normotensive | 0
appropriate fetal growth | 0
total weight gain of 14 pounds | 0
normal 20-week anatomy scan | 0
persistent productive cough | 0
shortness of breath | 0
intermittent nausea | 0
denied chest pain | 0
denied lower extremity swelling | 0
denied lower extremity pain | 0
tachycardia 111 beats per minute | 0
rupture of membranes | 0
closed cervix | 0
lungs clear to auscultation | 0
lower extremity edema 1+ | 0
urinary tract infection | 0
unknown GBS status | 0
started on steroid prophylaxis | 0
GBS prophylaxis | 0
ampicillin IV | 0
cefazolin | 0
cesarean section | 72
fever 40.2°C | 96
tachycardia | 96
suspicion of sepsis | 96
started on gentamicin | 96
started on clindamycin | 96
endometritis | 96
portable chest x-ray showed no acute cardiopulmonary disease | 96
blood cultures drawn | 96
blood cultures negative | 96
influenza tests negative | 96
RSV test negative | 96
urine Legionella antigen positive | 96
urine mycoplasma negative | 96
urine streptococcus antigen negative | 96
thyroid function tests normal | 96
lower extremity ultrasound negative for DVT | 96
transaminitis | 96
RUQ ultrasound normal liver | 96
common bile duct 0.5 cm | 96
questionable mild gallbladder wall thickening | 96
started on ceftriaxone | 96
started on azithromycin | 96
azithromycin changed to levofloxacin | 96
recurrent fever | 120
tachycardia up to 130 bpm | 120
transferred to ICU | 120
CT chest bilateral basilar infiltrates | 144
diagnosis of pneumonia | 144
ground glass opacity left upper lobe | 144
CT abdomen hepatic steatosis | 144
CT abdomen hepatomegaly | 144
ID consultation obtained | 144
switched to oral azithromycin | 168
treated with Zosyn for endometritis | 168
condition improved | 168
transferred out of ICU | 168
discharged | 216
complete additional 4 days of azithromycin | 216
blood pressure normal throughout | 216
transaminitis peaked on day 6 | 144
AST 813 U/L | 144
ALT 440 U/L | 144
INR normal | 144
bilirubin normal | 144
gastroenterology consultation | 144
serologic evaluation negative | 144
HSV-1 IgM positive | 216
HSV-2 IgM positive | 216
parvovirus B19 IgM positive | 216
ammonia normal | 144
repeat US hepatic steatosis | 144
hepatomegaly | 144
edema adjacent to gallbladder | 144
gallbladder normal | 144
common bile duct 2 mm | 144
hepatic arterial flow normal | 144
hepatic venous flow normal | 144
treated with NAC | 144
received loading dose | 144
received 15 follow-up doses | 144
refused last 2 doses | 144
Tylenol 2300 mg on day 4 | 96
refused transfer | 144
repeat LFT normalized | 216
LDH 212 U/L | 216
mild thrombocytopenia | 96
anemia | 96
nadired on postpartum day 1 | 96
nadired on day 3 | 144
haptoglobin normal | 144
LDH 615 U/L | 144
sodium 133 mEq/L | 144
