43 years old | 0
male | 0
myelodysplastic syndrome | 0
excess blasts-1 | 0
Kawasaki disease | -3960
hypertension | 0
hyperuricemia | 0
angina pectoris | 0
coronary artery lesions | -3960
surgery for coronary artery lesions | -3960
azacytidine | -72
COVID-19 IgG/IgM combined antibody test | 0
negative COVID-19 test | 0
PICC insertion | 0
local redness | 96
catheter removal | 96
broad-spectrum antimicrobial therapy | 96
piperacillin/tazobactam | 96
teicoplanin | 96
fever | 144
antimicrobials changed | 144
meropenem | 144
clindamycin | 144
right upper arm swelled | 144
difficulty bending elbow | 144
orthopedic surgeon consultation | 192
conservative treatment | 192
vital signs | 240
Glasgow Coma Scale | 240
temperature | 240
blood pressure | 240
heart rate | 240
respiratory rate | 240
oxygen saturation | 240
physical examination | 240
swelling and redness | 240
muscle pain | 240
tenderness | 240
blood investigations | 240
white blood cell count | 240
neutrophils | 240
hemoglobin | 240
platelet | 240
C-reactive protein | 240
total protein | 240
albumin | 240
aspartate aminotransferase | 240
alanine aminotransferase | 240
total bilirubin | 240
creatinine kinase | 240
blood urea nitrogen | 240
creatinine | 240
prothrombin time | 240
fibrinogen | 240
fibrin and fibrinogen degradation products | 240
D-dimer | 240
procalcitonin | 240
presepsin | 240
plain radiograph | 240
MRI | 240
necrotizing soft tissue infection | 240
septic shock | 240
urgent debridement surgery | 240
large fluid infusion | 240
noradrenaline infusion | 240
broad-spectrum antimicrobial agents | 240
meropenem | 240
daptomycin | 240
clindamycin | 240
posaconazole | 240
infectious myositis | 240
myonecrosis | 240
DVT of brachial vein | 240
catheter insertion site | 240
tissue culture | 240
histopathological examination | 240
muscle tissues | 240
surrounding exudate | 240
echo | 264
enhanced computed tomography | 264
thrombosis | 264
intravenous heparin | 264
ICU admission | 264
vital signs stable | 312
culture tests negative | 312
histopathological examination | 312
rehabilitation | 336
wound cleaning | 336
debridement | 336
negative-pressure wound therapy | 336
shoe-lace technique | 336
antimicrobials changed | 600
tosufloxacin | 600
posaconazole | 600
CRP levels negative | 840
wound closed | 1248
range of motion | 1814
elbow flexion | 1814
elbow extension | 1814