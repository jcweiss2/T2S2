Here is the extracted table of events with timestamps:

18 years old | 0
male | 0
Child–Pugh class C cirrhosis | 0
slipping on wet grass and falling on his left side | -4
admitted to the Emergency department | 0
glasgow coma score 15/15 | 0
vital signs within normal limits | 0
pulse rate 78/min | 0
RR 13/min | 0
BP 113/54 mm Hg | 0
SpO2 100% in air | 0
left hip tenderness | 0
no ecchymosis to the abdomen, flank or thigh | 0
radiograph of pelvis | 0
undisplaced fracture of his left acetabulum of both the anterior and posterior columns | 0
initial blood tests | 0
pH 7.271 | 0
base excess minus 7.3 | 0
PT 18.2 | 0
INR 1.5 | 0
APTT ratio 1.42 | 0
platelets 73 | 0
bilirubin 63 mmol/l | 0
Hb 124 g/l | 0
insertion of an 18 g intravenous cannula | 0
commenced warmed Hartmanns one litre infusion | 0
referred to the Orthopaedic on call team | 0
blood pressure dropped to 75/51 mm Hg | 0
tachycardic | 0
serum lactate was 9 mmol/l | 0
FAST examination | 0
intraabdominal fluid | 0
treated for sepsis | 0
intensive care, orthopaedic and general registrar attended the patient | 0
pH 7.227 | 0
base excess of −17.9 | 0
serum lactate of 16.3 mmol/l | 0
Hb 75 g/l | 0
arterial blood pressure was 90/60 mm Hg with a pulse rate 90/min | 0
left lower abdominal quadrant and upper thigh were now swollen with ecchymosis | 0
diagnosis of haemorrhaic shock | 0
massive transfusion pathway was activated | 0
four units of Blood | 0
four units of FFP | 0
two adult therapeutic doses of platelets | 0
ten units of cryoprecipitate | 0
noradrenaline infusion to maintain MAP > 65 mm Hg | 0
pelvic binder was in place but not tightened | 0
CT scan was deemed necessary | 0
on call radiology team and vascular surgeons were contacted | 0
CT abdomen confirmed the fracture of the left acetabulum | 0
significant haematoma on left pelvic sidewall adjacent to the fracture | 0
8 mm enhancing nodule suggestive of an internal iliac artery pseudoaneurysm | 0
ill-defined blush of contrast within the haematoma | 0
extra-peritoneal haematoma inseparable from the bladder | 0
cirrhotic liver | 0
incidental 6.7 cm infra-renal aortic aneurysm | 0
transferred to the intensive care unit | 0
CT Angiogram | 24
no arterial bleed | 24
prophylactic embolization | 24
gelfoam embolization of anterior and posterior division segmental branches of the left internal iliac artery | 48
10 lb skeletal traction was applied | 48
discharged to the orthopaedic ward | 120
uncontrollable bleeding from his pin site | 120
bleeding from his pin site while in skeletal traction | 120
removed and continuous pressure applied to the wound | 120
died on 30 January 2017 | 720