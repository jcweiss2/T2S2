79 years old | 0
woman | 0
presented to the Emergency Department | 0
slurred speech | 0
arm weakness | 0
deteriorating mobility | -2160
deteriorating cognition | -2160
deteriorating oral intake | -2160
not taking regular medications | 0
radioactive iodine treatment | -283104
hyperthyroidism | -283104
iatrogenic hypothyroidism | -283104
stopped levothyroxine | -126144
temperature 33.3°C | 0
heart rate 45 bpm | 0
blood pressure 170/99 mmHg | 0
oxygen saturations 90% | 0
GCS 9/15 | 0
dry flaky skin | 0
coarse hair | 0
frontal balding | 0
globally depressed reflexes | 0
hoarse voice | 0
peripheral oedema | 0
no palpable goitre | 0
CT head focal right cerebellar calcification | 0
no acute pathology | 0
stupor | 0
Na+ 127 mmol/l | 0
CRP 19 mg/l | 0
CK 586 IU/l | 0
TSH 51 mU/l | 0
T4 2.6 pmol/l | 0
T3 <0.8 pmol/l | 0
cortisol 1001 nmol/l | 0
re-warming | 0
broad-spectrum IV antibiotics | 0
possible aspiration pneumonia | 0
T4 25 μg NG route | 0
IV T3 10 μg three times a day | 0
regular hydrocortisone | 0
adrenal insufficiency | 0
no organ support | 0
critical care unit admission | 0
close monitoring | 0
treatment risks arrhythmia | 0
treatment risks myocardial infarction | 0
passed away | 672
recurrent hospital-acquired pneumonias | 672
NSTEMI | 672
per rectum bleed | 672
raised CK secondary to thyroid myositis | 672
myxoedema coma | 0
longstanding untreated hypothyroidism | 0
hypothermia | 0
infection | 0
stroke differential | 0
'cold' sepsis differential | 0
no consideration of thyroid dysfunction | 0
known hypothyroidism | 0
sepsis precipitating factor | 0
renal impairment | 0
hyponatremia | 0
hypoglycemia | 0
raised CK | 0
altered mental state | 0
precipitating event | 0
coarse dry hair | 0
alopecia | 0
dry skin | 0
generalized oedema | 0
macroglossia | 0
bradycardia | 0
delayed reflexes | 0
thyroid hormone replacement | 0
T4 replacement monotherapy | 0
T3 replacement | 0
IV T4 200–400 μg | 0
oral thyroxine | 0
constipation | 0
paralytic ileus | 0
combination treatment IV T3 | 0
NG T4 | 0
impaired T4-to-T3 conversion | 0
excess T3 cardiac side effects | 0
early improvement in neuropsychiatric symptoms | 0
IV T3 10–20 μg 8-hourly | 0
lower doses in elderly | 0
lower doses in ischemic heart disease | 0
hydrocortisone 50–100 mg IV | 0
coexistent adrenal insufficiency | 0
increased cortisol clearance | 0
multi-organ involvement | 0
critical care admission | 0
advanced age | 0
reduced consciousness level | 0
persistent hypothermia | 0
significant underlying precipitants | 0
myocardial infarction | 0
early treatment | 0
supportive measures | 0
infection treatment | 0
critical care environment | 0
