ingestion of two fresh tablets of Celphos (AlP) | -4
vomiting with 4–5 episodes | -4
pain in the abdomen | -4
agitated, anxious, and irritable | 0
pulse rate (PR) was not palpable | 0
blood pressure (BP) was not recordable | 0
heart rate (HR) was 110/minutes | 0
respiratory rate (RR) was 28/min | 0
oxygen saturation (SPO2) was 95% | 0
sinus tachycardia | 0
T wave inversion in lead 3 | 0
intravenous (IV) crystalloids | 0
IV magnesium sulphate 1 gm stat and 8 hourly | 0
IV calcium gluconate 8 hourly | 0
IV hydrocortisone 100 mg stat and 12 hourly | 0
IV dopamine | 0
noradrenaline | 0
gastric lavage with potassium permanganate (KMnO4) | 0
activated charcoal was kept in the stomach | 0
arterial blood gas (ABG) analysis showed a metabolic acidosis | 0
pH of 7.2 | 0
HCO3 of 8 mmol/L | 0
PCO2 of 33 mmol/L | 0
metabolic acidosis correction | 0
intubated | 0
shifted to an intensive care unit (ICU) | 0
BP was 60–80 mmHg (systolic) | 6
PR was 120/min | 6
RR was 20/min | 6
input/output was 3L/300 ml | 24
monomorphic ventricular tachycardia (VT) | 48
DC cardio-version of synchronised 150 J | 48
IV amiodarone 150 mg bolus and infusion | 48
normal sinus rhythm (NSR) | 48
cardiac bio-markers raised | 48
ABG showed a pH of 7.4 | 96
HCO3 of 18 mmol/L | 96
CO2 of 42 mmol/L | 96
BP was ranging from 70/50 mmHg to 90/60 mmHg | 96
blood urea was 100 mg/dl | 96
serum creatinine was 4.5 mg/dl | 96
urine output was 400 ml/24 hours | 96
aspartate amino-transferase/alanine amino-transferase (AST/ALT) was 80/90 IU/L | 96
alkaline phosphatase (ALP) was 200 U/L | 96
S bilirubin was 2.5 mg/dl | 96
liver and kidney involvement | 96
BP was 100/70 mmHg | 120
PR was 110/min | 120
RR was 22/min | 120
total leucocyte count (TLC) was 14000/mm3 | 120
polymorphonuclear leucocytosis | 120
Urea was 200 mg/dl | 120
S. creatinine was 7.5 mg/dl | 120
urine output was 400 ml/24 hours | 120
ABG showed re-appearance of acidosis | 120
pH was 7.1 | 120
HCO3 was 10 mmol/L | 120
haemodialysis | 120
haemodialysis | 168
blood urea after haemodialysis on the seventh day was 70 mg/dl | 168
creatinine was 4.0 mg/dl | 168
urine output improved to around 1200 ml/24 hours | 168
extubated | 144
shifted to a step down unit (SDU) | 192
vitals were normal | 192
liver and kidney functions were improving | 192
discharged | 336