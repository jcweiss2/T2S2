23 years old | 0
male | 0
admitted to the hospital | 0
fever | -120
highest temperature 39.1 °C | -120
received treatment at a local health clinic | -96
prescribed with cephalosporin antibiotics | -96
saw a doctor at Beijing Huairou District Hospital | -72
chest computed tomography (CT) scan | -72
large consolidation of the lower lobe of the right lung | -72
superior lobe of the left lung | -72
arterial blood gas analysis | -72
pH 7.476 | -72
PCO2 22 mmHg | -72
PO2 54.1 mmHg | -72
HCO3- 20.4 mmol/L | -72
FiO2 21% | -72
antigen of influenza A positive | -72
transferred to the general ICU | 0
history of atrial septal defect | -9360
history of ventricular septal defect | -9360
history of pulmonary artery stenosis | -9360
history of right ventricular double outlet | -9360
history of Tausing-Bing syndrome | -9360
modified Fontan operation | -9360
pulmonary orifice sutured | -9360
tricuspid valve sewn closed | -9360
left auricle connected with the pulmonary artery | -9360
recovered well after the operation | -9360
able to perform general physical activity | -9360
echocardiography at the regular visit | -1095
double outlet in the right ventricle | -1095
right atrial enlargement | -1095
aortic valve regurgitation | -1095
ejection fraction 50% | -1095
physical examination | 0
temperature 38.4 °C | 0
blood pressure 86/54 mmHg | 0
respiration rate 40 times/min | 0
pulse rate 110 times/min | 0
SPO2 80% | 0
breath sounds of both lungs thick and moist rales | 0
arrhythmia | 0
dropped-beat pulse | 0
respiratory failure | 0
septic shock | 0
skin wet, cold, and bluish | 0
laboratory examinations | 0
white blood cell count 11.89 × 10^9/L | 0
neutrophil percentage 84.94% | 0
hemoglobin 173.10 g/L | 0
hematocrit 48.70% | 0
platelet count 178.00 × 10^9/L | 0
sodium 128.5 mmol/L | 0
creatinine 279.6 µmol/L | 0
procalcitonin 4.51 ng/mL | 0
C-reactive protein 212.9 mg/L | 0
alanine aminotransferase 48.6 U/L | 0
aspartate aminotransferase 100.4 U/L | 0
total bilirubin 26.2 µmol/L | 0
direct bilirubin 21.4 µmol/L | 0
chest X-ray | 0
ventilator mode intermittent positive pressure ventilation | 0
FiO2 100% | 0
tidal volume 560 mL | 0
respiratory frequency 20 times/min | 0
positive end-expiratory pressure 10 cmH2O | 0
peak airway pressure 23 cm H2O | 0
moxifloxacin hydrochloride | 0
paramivir | 0
anti-infective drugs switched to cefoperazone-sulbactam sodium | 72
vancomycin hydrochloride | 72
voriconazole | 72
central venous pressure (CVP) 40 mmHg | 0
noradrenaline | 0
continuous renal replacement therapy | 0
protective lung ventilation strategy | 0
ventilation in prone position | 0
arterial blood gas analysis | 24
pH 7.193 | 24
PCO2 48 mmHg | 24
PO2 52 mmHg | 24
base excess -10 mmol/L | 24
lactate 1.34 mmol/L | 24
VV ECMO | 24
two vein indwelling catheters | 24
rotation speed 3100 turns/min | 24
blood flow volume 4.3 L/min | 24
oxygen flow volume 4.5 L/min | 24
FiO2 100% | 24
VV ECMO converted to VVA ECMO | 120
right femoral artery punctured and intubated | 120
combined deep venous catheters | 120
rotation speed 3800 turns/min | 120
blood flow volume 4 L/min | 120
oxygen flow volume 4 L/min | 120
FiO2 100% | 120
negative liquid equilibrium | 120
CVP decreased to 28 mmHg | 120
circulation tended to deteriorate | 120
noradrenaline dose adjusted | 120
cumulative positive balance 10000 mL | 168
CVP gradually increased to 35 mmHg | 168
noradrenaline dose tapered | 168
noradrenaline stopped | 336
oxygenator and circulation line replaced | 408
tracheotomy | 432
VVA ECMO equipment removed | 504
artificial ventilation withdrawn | 648
discharged from hospital | 720
follow-up | 1272