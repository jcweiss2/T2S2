70 years old | 0 | 0 
male | 0 | 0 
farmer | 0 | 0 
admitted to the hospital | 0 | 0 
high-grade fever | -120 | 0 
generalized body ache | -120 | 0 
headache | -120 | 0 
altered sensorium | -24 | 0 
joint pains | -120 | 0 
epigastric pain | -120 | 0 
no comorbidities | 0 | 0 
no drug addiction | 0 | 0 
no intoxication | 0 | 0 
inguinal lymphadenopathy | 0 | 0 
mild generalized rash | 0 | 0 
no eschar | 0 | 0 
hemodynamically stable | 0 | 0 
disoriented | 0 | 0 
no focal neurological deficit | 0 | 0 
no neck rigidity | 0 | 0 
acute febrile illness | 0 | 0 
undifferentiated fever | 0 | 0 
malaria test negative | 0 | 0 
dengue test negative | 0 | 0 
typhoid test negative | 0 | 0 
leptospira test negative | 0 | 0 
scrub typhus antigen card positive | 0 | 0 
scrub immunoglobulin M positive | 0 | 0 
diagnosis of scrub typhus | 0 | 0 
blood culture sterile | 0 | 0 
body fluid culture sterile | 0 | 0 
leukocytosis | 0 | 0 
mild hyperbilirubinemia | 0 | 0 
transaminitis | 0 | 0 
raised international normalized ratio | 0 | 0 
hepatitis B antigen negative | 0 | 0 
hepatitis C antibody negative | 0 | 0 
mild fatty infiltration of the liver | 0 | 0 
doxycycline treatment | 0 | 168 
defervescence | 48 | 48 
improved orientation | 48 | 48 
weakness of lower limbs | 96 | 96 
weakness progressed to upper limbs | 96 | 120 
absent deep tendon reflexes | 96 | 168 
flexor plantar responses | 96 | 168 
bladder incontinence | 96 | 168 
no bowel incontinence | 96 | 168 
breathing difficulty | 120 | 120 
respiratory distress | 120 | 120 
intubated | 120 | 120 
mechanical ventilation | 120 | 130 
MRI brain normal | 120 | 120 
MRI cervical spine normal | 120 | 120 
nerve conduction velocity test | 120 | 120 
motor sensory demyelinating polyneuropathy | 120 | 120 
Guillain-Barré syndrome diagnosis | 120 | 120 
cerebrospinal fluid analysis | 120 | 120 
intravenous immunoglobulin therapy | 120 | 125 
rifampicin treatment | 120 | 168 
improvement in weakness | 125 | 168 
improvement in respiratory parameters | 125 | 168 
weaned off ventilator | 130 | 130 
extubated | 130 | 130 
oral feeding started | 130 | 130 
limb physiotherapy | 130 | 168 
chest physiotherapy | 130 | 168 
shifted out of ICU | 168 | 168 
discharged from hospital | 168 | 168 
full neurological recovery | 168 | 168 
follow-up in outpatient department | 168 | 720 
no functional disability | 720 | 720