55 years old | 0
    farmer | 0
    admitted to a local county hospital | 0
    tick bite on left leg | -240
    fever | -168
    chills | -168
    obvious fatigue | -168
    body temperature normalized | -168
    fever repeatedly recurred within 48 hours | -120
    admitted to Lishui People's Hospital | 0
    temperature 40°C | -168
    respiratory rate 20 breaths/minute | -168
    blood pressure 116/65 mmHg | -168
    no ecchymosis or bleeding points in the skin | -168
    slightly coarse sounds in both lungs | -168
    no obvious dry and wet rales | -168
    heart rhythm regular | -168
    pain in the liver on percussion | -168
    palpable lymph node enlargement in the groin | -168
    total white blood cell count 3.1×10⁹/L | -168
    neutrophil count 2.48×10⁹/L | -168
    hemoglobin 138 g/L | -168
    platelet count 112×10⁹/L | -168
    C-reactive protein 66.7 mg/L | -168
    negative for hepatitis B surface antigen | -168
    normal urinalysis | -168
    chest CT revealed mild inflammation in both lungs | -168
    emphysema | -168
    sepsis | -168
    pneumonia | -168
    piperacillin 4.5 g every 8 hours for 2 days | -168
    no significant improvement | -168
    Tienam injection 1.0 every 8 hours for 2 days | -168
    no observable improvement | -168
    relapse | -72
    admitted to Department of Respiratory and Critical Care Medicine | 0
    temperature 38°C | 0
    pulse 67 beats/minute | 0
    blood pressure 113/69 mmHg | 0
    respiratory rate 21 breaths/minute | 0
    delirious | 0
    suspicious response to bending of neck | 0
    white blood cell count 3.5×10⁹/L | 0
    red blood cell count 4.38×10¹²/L | 0
    hemoglobin 132 g/L | 0
    platelet count 61×10⁹/L | 0
    erythrocyte sedimentation rate 17 mm/hour | 0
    prothrombin time 13.1 s | 0
    d-dimer 4546 µg/L | 0
    total protein 53.4 g/L | 0
    alanine aminotransferase 285 U/L | 0
    aspartate aminotransferase 235 U/L | 0
    total bile acids 30.9 µmol/L | 0
    C-reactive protein 130.8 mg/L | 0
    negative for blood plasmodia | 0
    negative for HIV | 0
    negative for hepatitis C | 0
    negative for anti-Epstein-Barr virus IgG | 0
    negative for syphilis | 0
    negative for pneumonia antibody | 0
    negative Widal test | 0
    negative Weil-Felix test | 0
    weakly positive urinary microalbumin | 0
    clear cerebrospinal fluid | 0
    weak positivity in Pandy's test | 0
    chloride 119 mmol/L | 0
    total protein 0.64 g/L | 0
    IgG 95 mg/dL | 0
    sterile cerebrospinal fluid culture | 0
    sterile blood culture | 0
    mild mitral valve reflux | 0
    tricuspid valve reflux | 0
    cardiac arrhythmia | 0
    calcification in left renal cortex | 0
    calcification in prostate | 0
    hepatomegaly | 0
    gallbladder wall thickening | 0
    abdominal cavity effusion | 0
    inflammation in both lungs | 0
    multiple small nodules in right and left lower lobes | 0
    patchy fibrosis in right middle lung lobe | 0
    patchy fibrosis in upper lobes of both lungs | 0
    emphysema | 0
    hepatomegaly | 0
    dilatation of intrahepatic lymphatic vessels | 0
    gallbladder wall edema | 0
    ascites | 0
    enlarged lymph nodes in abdominal cavity | 0
    enlarged lymph nodes in retroperitoneum | 0
    multiple low-density lesions in spleen | 0
    possible splenic infarction | 0
    small cysts in caudate hepatic lobes | 0
    small cyst in left kidney | 0
    calcification foci in prostate | 0
    bilateral pleural effusion | 0
    next-generation sequencing identified Coxiella burnetii | 168
    doxycycline hydrochloride enteric-coated capsules administered | 168
    compound glycyrrhizin injection | 168
    reduced glutathione injection | 168
    no fever | 264
    no chills | 264
    discharged | 264
    no side effects of therapy | 264
    doxycycline anti-infection sustained | 264
    compound glycyrrhizin/doxycycline treatment sustained | 264
    