78 years old | 0
woman | 0
diagnosed with hepatocellular carcinoma | 0
hypertension | 0
liver cirrhosis | 0
hepatitis C virus antibodies | 0
computed tomography revealed advanced HCC | 0
lenvatinib initiated at 8 mg/day | 0
treatment interrupted 2 months later | 720
proteinuria | 720
lenvatinib resumed at 4 mg/day | 7200
feeling unsteady on feet | -168
vomiting after ingesting small amounts of food | -168
presented with respiratory distress | -168
urge incontinence | -168
night sweats | -168
dehydration | 0
shock | 0
blood pressure not measurable | 0
heart rate 137 beats/min | 0
respiratory rate 33 breaths/min | 0
body temperature 36.4°C | 0
soft abdomen | 0
nontender abdomen | 0
no guarding | 0
white blood cells 15,700/μL | 0
hemoglobin 16.0 g/dL | 0
platelets 216,000/μL | 0
creatinine 2.90 mg/dL | 0
C-reactive protein 18.2 mg/L | 0
computed tomography showed free air bubbles | 0
emergency exploratory laparotomy | 24
peritonitis with purulent exudate | 24
focally necrotic perforation | 24
sigmoid colon perforation | 24
Hartmann's procedure | 24
sigmoid resection | 24
end colostomy | 24
transferred to intensive care unit | 24
died | 72
macroscopic examination of sigmoid colon | 24
histopathological examination | 24
infiltration of neutrophils | 24
hemorrhage around perforation site | 24
no malignant lesion | 24
lenvatinib-related bowel perforation suspected | 24
