41 years old | 0
male | 0
originally from West Africa | 0
questionable history of ventriculoseptal defect | 0
admitted to the hospital | 0
worsening exertional dyspnea | -336
palpitations | -336
loss of appetite | -336
lower extremity edema | -336
30 pounds weight loss | -336
temperature 98.8°F | 0
blood pressure 104/50 mm Hg | 0
heart rate 120/min | 0
respiratory rate 18/min | 0
oxygen saturation 98% | 0
chronically ill cachexic male | 0
BMI 21 kg/m2 | 0
jugular venous distension | 0
bilateral rales | 0
tachycardia | 0
RV heave | 0
4/6 pan-systolic murmur | 0
palpable thrill | 0
blood cultures obtained | 0
empiric intravenous antibiotics started | 0
transthoracic echocardiogram | 0
transesophageal echocardiogram | 0
large mass attached to aortic valve leaflet | 0
severe aortic regurgitation | 0
holodiastolic flow reversal in aorta | 0
mass attached to flail anterior mitral valve leaflet | 0
severe mitral regurgitation | 0
mass attached to pulmonic valve | 0
significant pulmonic regurgitation | 0
severe pulmonary hypertension | 0
Pulmonary Artery Systolic Pressure 65 mm Hg | 0
dilatation of aortic root | 0
fistula between aortic sinus and RV outflow tract | 0
blood culture revealed gram-positive cocci | 24
identified as Abiotrophia species | 24
transferred to tertiary care center | 24
right heart catheterization | 48
elevated filling pressures | 48
low cardiac index | 48
shunt fraction 2.1 | 48
emergent surgery | 72
aortic root abscess | 72
prophylactic grafting of left anterior descending coronary artery | 72
prophylactic grafting of obtuse marginal artery | 72
bio-prosthetic pulmonary valve replacement | 72
bio-prosthetic mitral valve replacement | 72
closure of congenital VSD | 72
closure of aorto-RV fistula | 72
aortic root replacement | 72
post-operative atrial fibrillation | 96
amiodarone therapy started | 96
intravenous penicillin | 0
intravenous gentamycin | 0
transesophageal echocardiogram post-intervention | 168
mild left ventricular dysfunction | 168
ejection fraction 45% | 168
competent bio-prosthetic valves | 168
repeat blood cultures negative | 168
discharged on intravenous vancomycin | 240