60 years old | 0
female | 0
bipolar affective disorder | 0
hypertension | 0
hypothyroidism | 0
paraplegia | 0
admitted to senior behavioral facility | -108
increasing confusion | -108
unable to communicate | -72
tachycardia | -72
tachypnea | -72
flushing | -72
diaphoresis | -72
fevers greater than 38°C | -72
transferred to Neurologic Critical Care Unit | 0
encephalopathic | 0
tachypneic | 0
tachycardic | 0
hypoxemic | 0
generalized rigidity | 0
2+/4 hyperreflexia | 0
leukocytosis | 0
acute kidney injury | 0
elevated serum creatinine phosphokinase | 0
procalcitonin elevated | 0
C-reactive protein levels within normal limits | 0
episodes of hypotension | 0
episodes of hypertension | 0
sepsis considered | 0
NMS considered | 0
serotonin syndrome considered | 0
non-convulsive status epilepticus considered | 0
other central nervous system pathology considered | 0
blood cultures obtained | 0
urine cultures obtained | 0
sputum cultures obtained | 0
lumbar puncture considered | 0
ziprasidone treatment | -168
haloperidol treatment | -168
lithium treatment | -168
duloxetine treatment | -168
oxybutynin treatment | -168
baclofen treatment | -168
IV bromocriptine treatment | 0
IV dantrolene treatment | 0
discontinuation of ziprasidone | 0
discontinuation of haloperidol | 0
discontinuation of lithium | 0
discontinuation of duloxetine | 0
discontinuation of oxybutynin | 0
cooling blanket | 0
antipyretics | 0
IV fluids | 0
electroencephalography | 12
generalized slowing | 12
no seizure activity | 12
magnetic resonance imaging | 12
no acute findings | 12
afebrile | 72
improved leukocytosis | 72
autonomic dysregulation resolved | 96
labile blood pressures ceased | 96
supplemental oxygen requirements ceased | 96
more awake | 96
less rigid | 96
dantrolene increased | 120
transferred out of NCCU | 120