35 years old | 0
female | 0
gave birth to healthy twins | 0
cesarean section | 0
threatened preterm delivery | -672
in vitro fertilization | -672
facial nerve paresis | -672
severe headache | 24
generalized tonic–clonic seizures | 24
loss of consciousness | 24
arterial blood pressure 195/110 mmHg | 24
heart rate 120 beats/min | 24
provisional diagnosis of eclampsia | 24
transferred to intensive care unit | 24
antihypertensive therapy | 24
intravenous infusion of magnesium sulphate | 24
ebrantil | 24
20% manitol | 24
diazepam | 24
bilateral vision loss | 48
complete blood count normal | 48
liver function tests normal | 48
clotting parameters normal | 48
electrocardiogram normal | 48
proteinuria 2+ | 48
ophthalmological examination | 48
cortical blindness | 48
mild right-sided facial nerve paresis | 48
multislice computed tomography scan | 48
hypodensity of posterior white matter | 48
vasogenic edema | 48
magnetic resonance imaging | 72
T2- and fluid-attenuated inversion recovery-weighted images | 72
hyperintense signals in white matter | 72
parietal and occipital regions | 72
junctions of vascular watershed zones | 72
antihypertensive medication | 72
enalapril maleate | 72
methyldopa | 72
human albumin | 72
follow-up ophthalmological examinations | 120
bilateral improvement of visual function | 120
best-corrected visual acuity 1.0 | 120
slit lamp examination normal | 120
fundus examination normal | 120
visual field image | 120
peripheral relative scotoma | 120
depressed sensitivity of paracentral left visual field | 120
follow-up magnetic resonance imaging | 168
regression of edema | 168
discrete residual changes | 168
posterior horns of side ventricles | 168
discharged from clinic | 216
oral antihypertensive therapy | 216
physical therapy for facial nerve paresis | 216