40 years old | 0
African-American | 0
female | 0
admitted to the emergency department | 0
history of chronic eczema | -720
previous alcohol abuse | -720
gout | -720
hypothyroidism | -720
worsening eruption | 0
intermittent diarrhea | 0
cutaneous eruption | -144
desquamation of the hands | -144
desquamation of the feet | -144
desquamation of the perioral skin | -144
desquamation of the perineal skin | -144
associated pain | -144
associated swelling | -144
hair loss | -144
increasing weakness | -576
fatigue | -576
unintentional weight loss | -576
70 pounds weight loss | -576
psychosocial habits | -720
1 to 2 glasses of wine a day | -720
smoking | -720
no significant family history | 0
not on any medications | 0
erythematous desquamative patches | 0
erosions | 0
crusted lesions | 0
diffuse nonscarring alopecia | 0
scaling patches on the vermillion lips | 0
punch biopsy of the left medial thigh | 0
psoriasiform epidermal spongiosis | 0
superficial perivascular lymphohistiocytic infiltrate | 0
diffuse hypogranulosis | 0
broad overlying parakeratosis | 0
ballooning degeneration of the spinous layer | 0
methicillin-resistant Staphylococcus aureus | 0
Escherichia coli sepsis | 0
pneumonia | 0
admitted to the intensive care unit | 0
ventilator respiratory support | 0
systemic antibiotics | 0
laboratory and imaging studies | 0
necrolytic acral erythema ruled out | 0
pellagra ruled out | 0
biotin deficiency ruled out | 0
low zinc levels | 0
antitransglutaminase antibodies positive | 0
antiendomysium antibodies positive | 0
diagnosis of celiac disease | 0
zinc deficiency | 0
gluten-free diet | 0
zinc sulfate | 0
resolution of gastrointestinal symptoms | 96
resolution of cutaneous symptoms | 96
discharged from the hospital | 96