60 years old | 0
male | 0
benign prostatic hyperplasia | 0
diabetes mellitus type 2 | 0
hemoglobin A1c of 7.8 | 0
history of urinary tract infections | 0
abdominal pain | -168
gross hematuria | -168
difficulty voiding | -168
worsening pain | -24
pneumaturia | -24
acute urinary retention | -24
tachycardia | 0
normotensive | 0
febrile to 102 °F | 0
rigors | 0
abdominal guarding | 0
rebound tenderness | 0
suprapubic tenderness | 0
lactic acid of 3.4 mMol/L | 0
white blood cell count of 7.9 K/μL | 0
hemoglobin of 8.9 g/dL | 0
serum sodium of 132 mEq/L | 0
creatinine of 2.27 mg/dL | 0
urinalysis demonstrated 11–50 WBC/hpf | 0
>100 RBC/hpf | 0
positive nitrates | 0
moderate leukocyte esterase | 0
free air under the diaphragm | 0
extensive pneumoperitoneum | 0
emphysematous cystitis | 0
bilateral hydronephrosis | 0
emphysematous pyelitis | 0
possible abscess near the dome of the bladder | 0
intravenous fluids administered | 0
broad-spectrum antibiotics administered | 0
exploratory laparotomy | 0
cystoscopy | 0
cloudy free fluid encountered | 0
culture of free fluid | 0
bladder perforation | 0
diffuse inflammation | 0
trabeculations | 0
diverticula | 0
partial cystectomy | 0
removal of necrotic bladder tissue | 0
abscess pockets | 0
bladder edges debrided | 0
suprapubic catheter placed | 0
urethral catheter placed | 0
bladder closed in two layers | 0
abdomen irrigated | 0
lactic acidosis resolved | 24
hemodynamically stable | 24
discharged | 96
trimethoprim-sulfamethoxazole prescribed | 96
failed voiding trials | 96
transurethral resection of the prostate scheduled | 96
urine culture grew Escherichia coli | 96
intra-abdominal culture grew Escherichia coli | 96
focal transmural necrosis | 96
acute and chronic inflammation | 96
intramural abscess | 96
serositis with fibrosis | 96