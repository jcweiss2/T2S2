18 years old | 0
male | 0
admitted to the hospital | 0
farmer | -672
atrial fibrillation | -672
benign prostatic hypertrophy | -672
trismus | -672
hypertonia | -672
C. tetani infection | -672
immunoglobulins | -672
tetanus vaccination | -672
metronidazole | -672
respiratory failure | -672
coma | -672
tracheostomy | -672
mechanical ventilation | -672
vasoactive support | -672
seizures | -672
baclofen | -672
midazolam | -672
diazepam | -672
electroencephalography | -672
ventilator-associated pneumonia | -672
Klebsiella pneumoniae | -672
methicillin-sensitive Staphylococcus aureus | -672
piperacillin-tazobactam | -672
worsening respiratory function | -672
opacity on chest radiography | -672
peripheral leukocytosis | -672
blood cultures | -672
tracheal secretion samples | -672
septic shock | -672
antibiotic therapy | -672
linezolid | -672
meropenem | -672
septic shock | -672
cholestasis | -672
acute edematous pancreatitis | -672
endoscopic treatment | -672
urinary tract infection | -672
multidrug-resistant organisms | -672
colistin | -672
amoxicillin-clavulanate | -672
tracheostomy closure | -672
pressure ulcers | -672
sarcopenia | -672
low handgrip strength | -672
appendicular skeletal mass | -672
Clostridioides difficile infection | -672
oral vancomycin | -672
atrial fibrillation with third-degree atrioventricular block | -672
single-chamber pacemaker implantation | -672
hyperkinetic delirium | -672
Pseudomonas aeruginosa bloodstream infection | -672
ceftazidime-avibactam | -672
amikacin | -672
SARS-CoV-2 | -672
remdesivir | -672
droplet isolation | -672
second recurrence of C. difficile | -672
fidaxomicin | -672
bloodstream infection | -672
Candida parapsilosis | -672
fluconazole-resistant | -672
MSSA | -672
Candida tropicalis | -672
caspofungin | -672
cefazolin | -672
bloodstream infection | -672
P. aeruginosa | -672
piperacillin-tazobactam | -672
aztreonam | -672
ceftazidime-avibactam | -672
cefepime | -672
tracheostomy closure | -672
nutritional supplementation | -672
malnutrition | -672
sarcopenia | -672
motor reconditioning | -672
postural transition | -672
aided transfers | -672
axial stability | -672
balance improvement exercises | -672
wheelchairs | -672
walkers | -672
rehabilitation | -672
ENT | -672
geriatric follow-up | -672
Clostridioides difficile infection | -672
oral vancomycin | -672
atrial fibrillation with third-degree atrioventricular block | -672
single-chamber pacemaker implantation | -672
hyperkinetic delirium | -672
Pseudomonas aeruginosa bloodstream infection | -672
ceftazidime-avibactam | -672
amikacin | -672
SARS-CoV-2 | -672
remdesivir | -672
droplet isolation | -672
second recurrence of C. difficile | -672
fidaxomicin | -672
bloodstream infection | -672
Candida parapsilosis | -672
fluconazole-resistant | -672
MSSA | -672
Candida tropicalis | -672
caspofungin | -672
cefazolin | -672
bloodstream infection | -672
P. aeruginosa | -672
piperacillin-tazobactam | -672
aztreonam | -672
ceftazidime-avibactam | -672
cefepime | -672
tracheostomy closure | -672
nutritional supplementation | -672
malnutrition | -672
sarcopenia | -672
motor reconditioning | -672
postural transition | -672
aided transfers | -672
axial stability | -672
balance improvement exercises | -672
wheelchairs | -672
walkers | -672
rehabilitation | -672
ENT | -672
geriatric follow-up | 0
diffuse erythematous or maculopapular eruption | 0
pruritus | 0
DRESS syndrome | 0
fever | 0
rash | 0
increased WBC count | 0
eosinophilia | 0
systemic involvement | 0
diffuse erythematous or maculopapular eruption | 0
pruritus | 0
DRESS syndrome | 0
fever persisted | 0
rash persisted | 0
discharged | 24