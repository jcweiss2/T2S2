17 years old | 0
male | 0
thorat pain | -168
odynophagia | -168
submitted for blood tests | -168
Hemoglobin: 7.0 g/dL | -168
Hematocrit: 21% | -168
WBC: 33 x 10^9 cells/L | -168
platelets: 38 x 10^9 cells/L | -168
Acute promyelocytic leukemia (M3) | -168
daunorubicin | -168
vesanoid | -168
extensive necrotic lesion | 0
unpleasant odor | 0
biopsy | 0
culture | 0
nonspecific chronic diffuse inflammation | 0
necrotic areas | 0
numerous bacteria | 0
Enterococcus spp | 0
Staphylococcus aureus | 0
Candida SP | 0
antibiotic therapy | 0
ceftazidime | 0
amicacin | 0
vancomycin | 0
fluconazole | 0
penicillin G | 0
pneumonia | 0
sepsis | 0
intensive care unit | 0
total recovery | 45
extensive loss of soft palate tissue | 45