Here is the table of events and timestamps:

35 years old | 0
pregnant | 0
34 + 4 wk past menstrual period | 0
fever | -10
cough | -10
aggravated dyspnoea | -5
positive urine pregnancy test | -40
natural conception | -40
conscious of foetal movement | -16
foetal movement | -16
fever with highest body temperature 39.2 ℃ | -10
cough | -10
yellow viscous sputum | -10
chest distress | -10
shortness of breath | -10
oral acetaminophen | -10
admitted to hospital | 0
body temperature 36.4 ℃ | 0
blood pressure 117/87 mmHg | 0
heart rate 130 beats/min | 0
respiratory rate 20 times/min | 0
cyanosis of the lip | 0
thick breathing sounds in both lungs | 0
right lower lung dry and wet rales | 0
regular heart rate | 0
no noises in the auscultation area of each valve | 0
gestational and symmetric abdominal type | 0
height 166 cm | 0
pre-pregnancy weight 46.5 kg | 0
body mass index 16.87 | 0
weight gain 8.8 kg during pregnancy | 0
uterine height 34 cm | 0
abdominal circumference 89 cm | 0
contractions sporadic and weak | 0
head presentation | 0
foetal heart sounds 142 beats/min | 0
intrapelvic and extrapelvic measurements normal | 0
pH 7.472 | 0
partial pressure of carbon dioxide 34.0 mmHg | 0
partial pressure of oxygen 56 mmHg | 0
sulfur dioxide 88.6% | 0
C-reactive protein (CRP) 186.33 mg/L | 0
erythrocyte sedimentation rate 69.00 mm/h | 0
procalcitonin (PCT) 2.24 ng/mL | 0
White blood cell (WBC) 18.29 × 10^9/L | 0
neutrophil % 90.10% | 0
lymphocyte 0.97 × 10^9/L | 0
Alkaline phosphatase 232 U/L | 0
total bilirubin 23.1 μmol/L | 0
albumin (ALB) 33.9 g/L | 0
K+ 2.93 mmol/L | 0
sodium 129 mmol/L | 0
chloride 89 mmol/L | 0
chest computed tomography (CT) multiple plaques, miliary foci, nodular foci with partial consolidation and cavities in the upper and lower lobes of both lungs | 0
obstetric ultrasound single viable foetus, head presentation, and oligohydramnios | 0
cardiac ultrasound and lower extremity vascular ultrasound no significant abnormalities | 0
first menarche at the age of 15 | -15
menstrual cycle regular, lasting for 3-4 d every 30 d | -40
last menstruation occurred on May 2, 2022 | -40
marriage at an appropriate age | -40
spouse healthy | -40
one pregnancy history, G2P1 | -40
full-term normal delivery of a female infant in 2006 | -40
Pregnancy combined with severe pneumonia novel coronavirus infection S. aureus infection type respiratory failure | 0
late pregnancy with 34 + 4 wk G2P1 left occiput anterior | 0
elderly second parturient women | 0
maternal lower weight | 0
oligohydramnion | 0
premature live baby | 0
electrolyte disturbance | 0
hypoproteinaemia | 0
cefoperazone sodium and sulbactam sodium for anti-infective therapy | 0
10 mg dexamethasone to promote foetal lung maturation | 0
oxyhemoglobin saturation continued to progressively decline | 0
foetal heart sounds 146 beats/min | 0
foetal distress | 0
dead foetus in the uterus | 0
caesarean section of the lower uterus | 0
mask oxygen inhalation to high-flow nasal cannula oxygen therapy | 0
fraction of inspired oxygen at 100% and a flow rate of 50 L/min | 0
cyanosis improved significantly | 0
oxyhemoglobin saturation increased to 95%-98% | 0
assisted ventilation by endotracheal intubation with a ventilator | 0
empirical antibiotic therapy to prevent infection by intravenous drip of meropenem and vancomycin | 0
symptomatic treatment of fluid and ALB infusion | 0
irrigation solution was collected and tested for metagenomic next-generation sequencing (mNGS) by bedside tracheoscopy | 0
S. aureus combined with novel coronavirus infection | 0
no acid-fast bacilli in the sputum tuberculosis smear | 0
tubercle bacillus-polymerase chain reaction (TB-PCR) and nontuberculosis mycobacterium-PCR were negative | 0
galactomannan experiments were normal | 0
continued intravenous drip of 1 g every 12 h (q12h) vancomycin and 1 g q8h meropenem | 0
anticoagulant therapy | 0
treatments to relieve the cough and reduce the amount of sputum | 0
nasal tube oxygen with a flow rate of 3-4 L/min | 24
chest CT showed multiple areas of inflammation in both lungs, mildly enlarged mediastinal lymph nodes and a small amount of bilateral pleural effusion | 24
CRP was 38.54 mg/L | 24
WBC count was 8.25 × 10^9/L | 24
PCT was 0.129 ng/mL | 24
potassium was 4.04 mmol/L | 24
D-dimer was 2.44 mg/L | 24
TB-PCR was negative | 24
antibiotics were adjusted to sitafloxacin 50 mg twice daily | 48
patients’ condition was stable | 72
discharged from the hospital without special treatment | 72