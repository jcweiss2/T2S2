54 years old | 0
male | 0
smoking | 0
hypothyroidism | 0
T2N2bM0 squamous cell carcinoma | 0
human papillomavirus positive | 0
metastases to the cervical lymph nodes | 0
enrolled in the OPTIMA trial | 0
carboplatin/abraxane induction chemotherapy | -168
good imaging response | -168
complete resolution of primary tongue tumor | -168
decrease in size of cervical lymph nodes | -168
minimal side effects from chemotherapy | -168
admitted for inpatient chemoradiotherapy | 0
5-FU | 0
paclitaxel | 0
hydroxyurea | 0
fever | 24
pancytopenia | 24
intractable diarrhea | 48
vomiting | 48
hydroxyurea dose-decreased | 48
hydroxyurea held | 72
septic shock | 96
progressive desquamative skin lesions | 96
acute kidney failure | 96
sustained pancytopenia | 96
transferred to intensive care unit | 120
intubated | 120
transitioned to comfort care | 120
expired | 192
autopsy performed | 192
skin lesions | 192
toxic epidermal necrolysis | 192
bone marrow examination | 192
markedly hypocellular bone marrow | 192
diminished trilineage hematopoiesis | 192
virtually no megakaryocytes | 192
diffuse acute tubular necrosis | 192
gastrointestinal tract severely damaged | 192
post-mortem blood cultures positive for Stenotrophomonas maltophilia | 192
bilateral lung cultures positive for Stenotrophomonas maltophilia | 192
DNA analysis by next generation sequencing | 192
DPYD*2A/c.1905+1G>A mutation | 192
homozygous for nonfunctional alleles | 192
DPD deficiency | 192