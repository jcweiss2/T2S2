19 years old | 0
    male | 0
    admitted to a toxicology ward | 0
    significant sleepiness | 0
    unclear speech | 0
    drinking bout lasting 3 months | -2160
    alcohol addiction for 5 years | -43800
    Tourette syndrome | -43800
    clinical symptoms of pneumonia | -2160
    rapid deterioration of general condition | -2160
    required intubation | -2160
    mechanical ventilation | -2160
    echocardiographic examination revealed vegetations on heart valves | -2160
    transferred to intensive care unit | -2160
    intubated | -2160
    mechanically ventilated | -2160
    sedated with midazolamum | -2160
    sedated with fentanyl | -2160
    transthoracic echocardiography (TTE) | -2160
    grade 4 mitral insufficiency | -2160
    vegetation 1.2 × 1.6 cm on anterior cusp | -2160
    rupture of tendinous cords of anterior cusp | -2160
    vegetation 1.0 cm on posterior cusp | -2160
    aortic valve cusps marginal thickening | -2160
    vegetation on aortic valve | -2160
    grade 1 aortic insufficiency | -2160
    tricuspid valve insufficiency | -2160
    grade 1 central regurgitation jet | -2160
    suspected vegetation on tricuspid valve | -2160
    empiric antibiotic therapy (imipenem, vancomycin, clindamycinum) | -2160
    bacteriological analysis of venous blood | -2160
    bacteriological analysis of urine | -2160
    bacteriological analysis of bronchial secretions | -2160
    sterile cultures | -2160
    dental consultation | -2160
    numerous inflammatory foci in oral cavity | -2160
    extraction of 8 carious teeth | -2160
    7 days of antibiotic therapy | -2160
    presence of mobile vegetations on valves | -2160
    risk of embolization | -2160
    transferred to operating room | -2160
    surgical procedure using extracorporeal circulation (ECC) | -2160
    median sternotomy | -2160
    ascending aorta cannulated | -2160
    venous cannulas placed in caval veins | -2160
    aortic cross-clamping | -2160
    administration of crystalloid cardioplegic solution | -2160
    right ventricle opened | -2160
    tricuspid valve removed | -2160
    interatrial septum incised | -2160
    bicuspid valve removed | -2160
    aortic valve removed through aorta incision | -2160
    valve dysfunction (insufficiency, cusp perforation, vegetation) | -2160
    implantation of bioprostheses: Medtronic Hancock II Porcine 29 (mitral), Edwards Lifesciences C-E Perimount 21 (aortic), Medtronic Hancock II Porcine 33 (tricuspid) | -2160
    aortic cross-clamping time 161 minutes | -2160
    ECC time 224 minutes | -2160
    total surgery time 340 minutes | -2160
    transferred to recovery room | -2160
    hemodynamically stable | -2160
    requiring moderate catecholamines | -2160
    third postoperative day | -72
    mediastinal drains removed | -72
    intubated | -72
    mechanically ventilated | -72
    transferred to intensive care unit | -72
    antibiotic therapy continued | -72
    cultures from blood sterile | -72
    cultures from valves sterile | -72
    14th day of ICU stay | 336
    extubated | 336
    23rd postoperative day | 552
    general condition deteriorated | 552
    high fever | 552
    transferred to cardiology ward | 552
    sepsis diagnosed | 552
    bacteriological tests | 552
    Pseudomonas aeruginosa cultured from central venous catheter tip | 552
    Pseudomonas aeruginosa cultured from urine | 552
    Pseudomonas aeruginosa cultured from bronchial secretions | 552
    Pseudomonas aeruginosa cultured from peripheral venous blood | 552
    targeted antibiotic therapy (imipenem, Brulamycin) | 552
    no clinical improvement | 552
    fever persisted | 552
    weakness persisted | 552
    transesophageal echocardiography (TEE) | 552
    vegetation on aortic valve bioprosthesis | 552
    computed tomography (CT) of chest, head, abdomen | 552
    X-ray of chest | 552
    no inflammatory lesions | 552
    no metastatic abscesses | 552
    echocardiographic examination | 552
    cardiac surgical consultations | 552
    decision to replace aortic valve bioprosthesis | 552
    46th day after initial surgery | 1104
    transferred to operating room | 1104
    connected to ECC | 1104
    aortic cross-clamping | 1104
    administration of cardioplegia | 1104
    right atrium opened | 1104
    interatrial septum opened | 1104
    mitral bioprosthesis checked | 1104
    tricuspid bioprosthesis checked | 1104
    no vegetation found | 1104
    aorta opened | 1104
    conglomerate of vegetation on non-coronary cusp | 1104
    aortic valve bioprosthesis removed | 1104
    Edwards Lifesciences C-E Perimount 21 reimplanted | 1104
    aortic cross-clamping time 92 minutes | 1104
    ECC time 140 minutes | 1104
    transferred to recovery room | 1104
    extubated after 19 hours | 1133
    antibiotic therapy continued | 1133
    Pseudomonas aeruginosa cultured from removed aortic valve bioprosthesis | 1133
    postoperative blood cultures sterile | 1133
    12th day after reoperation | 1536
    transferred to cardiac rehabilitation hospital | 1536
    oral anticoagulation recommended for 3 months | 1536
    antibiotic therapy continued | 1536
    control echocardiographic examination on 30th day | 1680
    normal function of all bioprostheses | 1680