31 years old | 0
male | 0
admitted to the hospital | 0
high fever | 0
sore throat | 0
previously healthy | 0
no medications | 0
lived with wife and 11-month-old baby boy | 0
kept a dog | -744
son had high fever | -1344
son had strawberry tongue | -1344
son had desquamation of fingertips | -1344
son's symptoms resolved | -1344
body temperature elevated to 39℃ | 0
swollen and reddened pharynx | 0
erythema of trunk and right thigh | 0
negative streptococcal antibody tests | 0
ampicillin/sulbactam administered | 0
septic shock | 0
noradrenalin support | 0
referred to hospital | 0
no gastrointestinal symptoms | 0
well oriented | 0
blood pressure 112/54 mmHg | 0
heart rate 110 beats/min | 0
respiratory rate 24 breaths/min | 0
oxygen saturation 96% | 0
body temperature 37.3℃ | 0
conjunctivae congested | 0
erythema on right lower limb | 0
increased white blood cell count | 0
elevated erythrocyte sedimentation rate | 0
elevated C-reactive protein | 0
elevated total and direct bilirubin | 0
elevated serum ferritin | 0
elevated soluble interleukin-2 receptor | 0
elevated brain natriuretic peptide | 0
elevated procalcitonin | 0
decreased serum total protein | 0
decreased serum albumin | 0
normal platelet count | 0
blood urine and cerebrospinal fluid cultures unremarkable | 0
contrast-enhanced CT scanning | 0
bilaterally enlarged posterior cervical lymph nodes | 0
pulmonary congestion | 0
mild splenomegaly | 0
no lymphadenopathy | 0
treatment initiated for septic shock | 0
IV meropenem and gamma-globulin administered | 0
antibiotic changed to levofloxacin and clindamycin | 48
fever not resolved | 48
minocycline added | 120
fever and general condition improved | 120
moved to general ward | 216
bilateral desquamation of fingertips | 216
met clinical criteria for Kawasaki disease | 216
increasing platelet count | 216
coronary CT angiography | 384
no lesions | 384
cardiac ultrasonography | 1440
unremarkable | 1440
paired serum samples negative for anti-leptospiral antibodies | 72
discharged | 480
no signs of recurrence | 480
streptococcal or staphylococcal toxic shock syndromes considered | 0
did not meet criteria for toxic shock syndromes | 0
increase in platelet count during recovery | 216
FESLF suspected | 216
paired serum samples negative for anti-YPM antibodies | 72
agglutination reaction test positive for Y. pseudotuberculosis antibody | 96
diagnosed with FESLF | 216
son had similar symptoms | -1344
domestic transmission suspected | 0
contaminated well water possible source | 0
dog possible source | 0
refractory shock possibly due to YPM | 0
YPM has superantigen activity | 0
negative result for anti-YPM antibodies possibly false-negative | 72
treatment not established | 0
Y. pseudotuberculosis susceptible to antibiotics | 0
third-generation cephalosporins or fluoroquinolones recommended | 0
treatment recommended for 3 weeks | 0