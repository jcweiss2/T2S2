44 years old | 0
male | 0
hypertension | 0
chronic glomerulonephritis | 0
stage III chronic kidney disease | 0
stable eGFR of 30-35 | 0
amlodipine | 0
doxazosin | 0
ramipril | 0
presented to the emergency department | 0
shortness of breath | 0
loose stools | 0
fatigue | 0
hypoxia | 0
oxygen saturations 84% on air | 0
febrile (39.4°C) | 0
dyspnoeic | 0
respiratory rate 33/min | 0
placed on 15L oxygen therapy | 0
septic screen performed | 0
intravenous antibiotics | 0
fluids given | 0
urinary output monitoring | 0
chest radiographs patchy consolidation left lung base | 0
oxygen saturation 92% on 15L oxygen | 0
deteriorating work of breathing | 0
sedation | 0
intubation | 0
ventilation | 0
transferred to ICU | 0
remained sedated | 0
ventilated for 11 days | 264
repeat chest radiograph progression pulmonary opacification | 264
oxygen requirement peaked at day 4 | 96
hypoxaemia improvement | 96
slow weaning commenced | 96
respiratory viral PCR positive SARS-CoV-2 | 0
negative adenovirus | 0
negative influenza A | 0
negative influenza B | 0
negative parainfluenza viruses | 0
negative rhinovirus | 0
negative human enterovirus | 0
negative urinary pneumococcal antigen | 0
negative legionella antigen testing | 0
negative blood-borne virus | 0
negative sickle cell screening | 0
successfully extubated | 264
slow wean off oxygen therapy to room air | 264
recovery with regular physiotherapy | 264
post-extubation chest radiograph residual patches airspace opacification | 264
discharged | 264
persistent exercise limiting dyspnoea | 264
unable to return to functional baseline for 5 months | 264
developed malaise | 264
odynophagia | 264
after 2 weeks developed anterior neck swelling | 528
persisting pain | 528
no intervening illness | 528
10-day course oral penicillin antibiotics | 528
presented again with painful goitre | 528
pain on swallowing | 528
no signs of infection | 528
pain initially right side | 528
pain moved to contralateral side | 528
thyrotoxicosis | 528
slight weight loss | 528
general malaise | 528
mild autonomic symptoms of heat intolerance | 528
no tremor | 528
no palpitations | 528
no anxiety | 528
increased resting heart rate 90 bpm | 528
hyperthyroid biochemical picture | 528
antithyroid peroxidase antibodies positive | 528
raised inflammatory markers | 528
prescribed propranolol 40 mg once daily | 528
follow-up thyroid function testing | 528
ultrasound imaging of the neck | 528
geographic hypoechoic areas thyroid lobes | 528
minimal colour flow Doppler signal | 528
reactive cervical lymph nodes | 528
normal salivary glands | 528
commenced on propranolol | 528
simple analgesia | 528
paracetamol | 528
nonsteroidal anti-inflammatory drug (ibuprofen) | 528
hyperthyroid biochemical picture persisted at 3 weeks | 528
TSH 0.006 mIU/L | 528
free T4 21.7 pmol/L | 528
free T3 5.2 pmol/L | 528
anterior neck pain settled after 6 weeks | 528
swelling reduced | 528
pain reduced | 528
symptoms of thyrotoxicosis improved | 528
resolution of general malaise | 528
resolution of hot flushes | 528
corticosteroids not used | 528
antithyroid medications not used | 528
repeat TSH at 8 weeks | 1344
mild hypothyroid biochemical picture | 1344
hypothyroid period lasted 4 weeks | 1344
normalisation of thyroid hormones | 1344
serum TSH concentration on day 2 of intubation | 48
TSH 1.4 mIU/L | 48
onset of subacute thyroiditis after clinical resolution of SARS-CoV-2 | 528
negative SARS-CoV-1 hypothyroidism reports | 528
written informed consent | 528
no conflicts of interest | 528
no funding received | 528
