61 years old | 0
African-Canadian | 0
female | 0
admitted to the hospital | 0
fever | 0
dyspnea | 0
pneumonia | 0
chronic kidney disease | -672
previous pyoderma gangrenosum | -672
left above-knee amputation | -672
diabetes mellitus | -672
hypertension | -672
osteoarthritis | -672
sarcoidosis | -672
permanent hemodialysis catheter inserted | -168
hemodialysis started | -168
discharged | -168
diarrhea | -168
vomiting | -168
blood pressure 157/79 mm Hg | 0
heart rate 97 beats per minute | 0
respiratory rate 20 breaths per minute | 0
temperature 38.3°C | 0
oxygen saturation 98% | 0
purulent discharge around catheter exit site | 0
redness around catheter exit site | 0
induration along the tunnel | 0
tenderness along the tunnel | 0
admitted with diagnosis of dialysis catheter tunnel infection | 0
intravenous cloxacillin 2 g every 6 hours | 0
vancomycin 15 mg/kg bolus | 0
catheter removed | 0
catheter tip sent for culture | 0
high-grade fever | 24
leukocytosis | 24
swelling at catheter tunnel exit site expanded | 24
ulcerated with multiple points of purulent discharge | 24
new painful nodular lesion on abdominal wall | 48
ulcerated | 48
blood cultures repeated | 48
sterile cultures | 48
broadened antibiotic coverage to piperacillin/tazobactam | 72
diagnosis of pyoderma gangrenosum entertained | 168
consultation with rheumatology | 168
decision to avoid biopsy | 168
diuretics maximized | 168
stable without dialysis for 11 days | 168
initiation of steroids for pyoderma delayed | 168
hemodynamic instability | 192
BP 94/39 mm Hg | 192
acute alteration of mental status | 192
C-reactive protein 335 mg/L | 192
leukocyte count 28.7 × 10^9/L | 192
normal serum lactate | 192
resuscitated with intravenous fluids | 192
transferred to intensive care unit | 192
computed tomography of chest, abdomen, and pelvis | 192
left lower lobe consolidation | 192
mediastinal lymphadenopathy | 192
intravenous hydrocortisone 50 mg every 6 hours | 192
antibiotics continued unchanged | 192
fever resolved | 216
pain at site of lesions improved | 216
new tunneled dialysis line inserted | 216
hemodialysis resumed | 216
intravenous hydrocortisone changed to oral prednisone 50 mg/day | 216
piperacillin/tazobactam stopped | 216
intravenous vancomycin continued for 4 weeks | 216
discharged | 672
skin ulceration continued to improve | 1344
ulcers almost completely healed | 1344