53 years old| 0
male | 0
hypertension | 0
hypercholesterolemia | 0
bioprosthetic aortic valve replacement | 0
bicuspid aortic valve | 0
acute abdominal pain | -4320
lower extremity pain | -4320
weakness | -4320
right neck pain | -4320
low-grade fevers | -1440
sweats | -1440
malaise | -1440
dysphagia | -1440
febrile | 0
bilateral cold lower extremities | 0
absent femoral pulses | 0
ascending aortic pseudoaneurysm | 0
embolic occlusions | 0
prosthetic aortic valve | 0
intravenous vancomycin | 0
cefepime | 0
limb ischemia | 0
emergency laparotomy | 24
surgical thrombectomies | 24
bilateral lower limb fasciotomies | 24
mechanical ventilation | 24
vasopressors | 24
renal replacement therapy | 24
multiple acute infarcts | 24
intraparenchymal hemorrhages | 24
subarachnoid hemorrhages | 24
infiltrates with pigmented septate fungal hyphae | 30
melanin in the fungal cell wall | 30
broad-spectrum antifungal therapy | 30
liposomal amphotericin B | 30
intravenous voriconazole | 30
intravenous micafungin | 30
negative bacterial cultures | 30
negative fungal cultures | 30
Karius test | 30
Curvularia species detected | 30
fungal culture growth | 30
Curvularia alcornii identification | 30
ascending aorta replacement | 504
hemi-arch replacement graft | 504
biological Bentall aortic root and valve replacement | 504
large mycotic aneurysm | 504
fungal balls | 504
amphotericin B susceptibility | 504
voriconazole susceptibility | 504
fluconazole susceptibility | 504
itraconazole susceptibility | 504
ketoconazole susceptibility | 504
right neck swelling | 1440
increased pulsatility | 1440
right external carotid artery pseudoaneurysm | 1440
open right external carotid artery ligation | 1992
septate hyphae | 1992
liposomal amphotericin B completion | 1992
micafungin completion | 1992
suppressive oral voriconazole | 1992
progressive left leg pain | 2448
left leg numbness | 2448
fever | 2448
voriconazole level | 2448
bilateral iliac artery pseudoaneurysms | 2448
bilateral iliac artery coil embolization | 2448
liposomal amphotericin B restart | 2448
micafungin restart | 2448
posaconazole | 2448
arterial pseudoaneurysms | 2448
emboli | 2448
persistent fever | 2448
comfort care | 3600
death | 3600
