69 years old | 0
male | 0
Chinese | 0
admitted to the hospital | 0
hypertension | -672
coronary artery disease | -672
stage 4 chronic kidney disease | -672
diarrheal illness | -168
no fever | -168
no nausea | -168
no abdominal pain | -168
no jaundice | -168
septic shock | 12
transferred to the Medical Intensive Care Unit | 12
intravenous ceftriaxone | 12
blood cultures returned positive for P. aeruginosa | 24
meropenem | 24
sharply defined erythematous plaques | 48
erythematous plaques spread | 48
tense bullae | 60
bullae containing serous fluid | 60
bullous drug reaction | 48
bullous erysipelas | 48
septic vasculitis | 48
biopsy | 60
histological examination | 72
partial necrosis of the epidermis | 72
sub-epidermal blistering | 72
microthrombi | 72
neutrophilic infiltrate | 72
nuclear dust | 72
Gram-negative bacilli | 72
fluid culture of a needle aspirate | 72
P. aeruginosa | 72
aggressive fluid resuscitation | 72
high vasopressor support | 72
appropriate antibiotic therapy | 72
severe sepsis | 96
ST elevation myocardial infarction | 120
disseminated intravascular coagulopathy | 168
intracranial bleeding | 168
death | 168