65 years old | 0
female | 0
admitted to the oncology clinic | 0
abdominal pain | -30
pancreatic head lesion | -30
history of stage IIIA lung cancer | -810
smoking history | -810
hypertension | -810
hypothyroidism | -810
dyslipidemia | -810
spiculated suprahilar 4.5 × 2.6 cm right upper lobe (RUL) nodule | -810
multiple sub-centimeter left lung nodules | -810
augmented activity in the RUL mass | -810
NSCLC | -810
adenocarcinoma | -810
program death ligand-1 expression 15% | -810
carboplatin | -630
paclitaxel | -630
radiation therapy | -630
decrease in the RUL mass | -420
adjuvant immunotherapy with durvalumab | -420
pneumonitis | -390
steroid taper | -390
increase in the RUL mass | -270
increase in the RUL mass | -180
abdominal and pelvic CT scan | -30
mass in the head of the pancreas | -30
pancreatic ductal dilatation | -30
endoscopic ultra-sound-guided biopsy of the pancreatic head mass | 0
tumor cells with nuclear pleomorphism | 0
CK7 positivity | 0
TTF-1 positivity | 0
Napsin-A positivity | 0
CDX-2 negativity | 0
KOC negativity | 0
synaptophysin negativity | 0
Smad-4 mixed staining pattern | 0
lung adenocarcinoma metastasized to the pancreas | 0
AST 35 U/L | 0
ALT 23 U/L | 0
ALP 74 U/L | 0
total bilirubin 0.5 mg/dL | 0
direct bilirubin 0.2 mg/dL | 0
CA 19.9 22.5 U/mL | 0
PET/CT scan | 30
fluorodeoxyglucose-avid mass in the pancreatic head | 30
increased uptake in the porta hepatis | 30
brain MRI scan | 30
palliative radiation therapy | 90
combination chemotherapy with carboplatin and pemetrexed | 90
generalized weakness | 120
dyspnea at rest | 120
electrolyte derangements | 120
acute anemia | 120
hemoglobin nadir of 6.9 g/dL | 120
transfusion | 120
new 9 mm left lower lobe nodule | 120
staging PET/CT scan | 210
decreased metabolic activity in the pancreatic mass | 210
metabolic activity in the new left lower lobe nodule | 210
fatigue | 210
rapid response | 240
saturating at 87% on 3 L of oxygen via nasal cannula | 240
accessory muscles | 240
blood pressure of 84/70 | 240
heart rate of 138 | 240
increased dyspnea | 240
cough | 240
generalized weakness | 240
right lung consolidation | 240
loculated pleural effusion | 240
treatment for acute hypoxic respiratory failure | 240
sepsis secondary to pneumonia | 240
broad-spectrum antibiotics | 240
oxygen supplementation | 240
bilevel-positive airway pressure | 240
episode of altered mentation | 246
worsening hypoxemia | 246
vasopressor support | 246
palliative medicine team | 246
inpatient hospice care | 246
death | 252