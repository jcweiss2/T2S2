77 years old | 0  
    male | 0  
    hypertension | 0  
    diabetes | 0  
    ischemic heart disease | 0  
    captopril 25 mg tablet twice daily | 0  
    metformin 500 mg tablet twice daily | 0  
    aspirin 100 mg tablet once daily | 0  
    atorvastatin 20 mg tablet | 0  
    admitted to the emergency department | 0  
    progressive weakness in lower limbs | -72  
    retention of urine | -72  
    loss of all sensations in lower limbs up to umbilicus level | -72  
    febrile illness | -168  
    no shortness of breath | -168  
    no cough | -168  
    general examination | 0  
    full consciousness | 0  
    wakeful | 0  
    alert | 0  
    normal vital signs | 0  
    low-grade fever (38°C) | 0  
    no dyspnea | 0  
    no tachypnea | 0  
    chest auscultation fine crackles | 0  
    normal S1 heart sounds | 0  
    normal S2 heart sounds | 0  
    abdomen soft | 0  
    palpable distended bladder | 0  
    neurological examination | 0  
    normal higher cerebral function | 0  
    normal speech | 0  
    intact cranial nerves | 0  
    upper limb normal strength (5/5) | 0  
    reflexes +2 | 0  
    normal sensory examination | 0  
    lower limb flaccid paralysis (0/5) | 0  
    hypotonia | 0  
    reflexes grade 0 | 0  
    bilateral mute planter reflex | 0  
    extensor reflexes after 2 days | 48  
    sensory level at T10 | 0  
    loss of all sensations below T10 | 0  
    retention of urine | 0  
    elevated WBC count | 0  
    lymphopenia | 0  
    elevated renal indices | 0  
    chest CT showing COVID-19 features | 0  
    cervical dorsal MRI normal | 0  
    lumbosacral spine MRI normal | 0  
    negative PCR for CMV | 0  
    negative PCR for EBV | 0  
    negative PCR for HSV-1 | 0  
    negative PCR for HSV-2 | 0  
    negative serology for HCV | 0  
    negative serology for Mycoplasma pneumoniae | 0  
    negative serology for Brucella | 0  
    negative Quanti FERON-TB Gold test | 0  
    isolation | 0  
    methylprednisolone 1 g i.v. | 0  
    insulin therapy | 0  
    ceftriaxone 1 g i.v. | 0  
    azithromycin 250 mg capsules | 0  
    referral to COVID-19 hospital | 24  
    positive SARS-CoV-2 RT-PCR | 24  
    progressive deterioration | 48  
    shortening of breath | 48  
    admitted to ICU | 48  
    mechanical ventilation | 48  
    death | 96  
    multiorgan failure | 96  
    septicemia | 96  
    Babinski signs | 48  
    inflammatory myelopathy | 0  
    respiratory failure | 96  
    