25 years old | 0
male | 0
penetrating sharp injury with nail to left heel | -480
lockjaw | -288
muscle spasms in left lower extremity | -288
vaccination history negative | 0
awake | 0
trismus | 0
opisthotonos | 0
generalized attacks every 3-4 minutes in left leg | 0
injection of human anti-tetanus immunoglobulin (Hyper-Tet 250 U) | 0
injection of tetanus-diphtheria toxoid | 0
admitted to ICU | 0
midazolam infusion | 0
morphine infusion | 0
feeding via nasogastric tube | 0
severe spasms | 0
risk of rhabdomyolysis | 0
hydration with half saline 4 L/day | 0
bicarbonate infusion | 0
metronidazole 500 mg/qid/iv | 0
temperature 38°C | 72
tazocine 3.375 g/qid | 72
ciprofloxacin 500 mg iv | 0
positive urine culture (Escherichia coli > 100,000) | 0
severe generalized spasm | 0
pain | 0
intubated | 0
pancronium 4 mg loading dose | 0
pancronium 2 mg/hour | 0
percutaneous dilatational tracheostomy | 240
muscle relaxant discontinued | 360
spastic attacks in left leg continued | 360
high doses of sedative agents | 360
ventilation and oxygenation disrupted | 360
unable to extubate | 360
baclofen prescribed | 360
ultrasound-guided sciatic nerve block | 432
pain score decreased to less than 2 | 432
pain relieved | 432
extubated | 432
tachycardia | 0
stable blood pressure | 0
normal routine laboratory data | 0
normal liver function test | 0
creatine phosphokinase raised to 4500 IU/L | 0
left ICU with good general condition | 432
no consciousness impairment | 0
no dysphagia | 0
no laryngospasm | 0
no spasm of respiratory tract muscles | 0
no cardiorespiratory arrest | 0
gag intact before intubation | 0
fed by tube | 0
spastic attacks continued | 360
intermittent low dose of midazolam | 432
analgesia continued for 48 hours | 432
pain tolerable after nerve block relief | 480
no need for opioid-analgesic agents | 480
