15 months old | 0
male | 0
admitted to the hospital | 0
Wiskott–Aldrich syndrome | -672
thrombocytopenia | -672
genetic studies | -672
four-base-pair deletion in intron-8 | -672
no protein expression of WAS | -672
unaffected sister was not a human leukocyte antigen match | -672
required platelets transfusions | -336
worsening petechiae | -336
intermittent hematochezia | -336
intravenous immunoglobulin therapy | -336
prophylactic trimethoprim-sulfamethoxazole | -336
admitted for preconditioning therapy | -24
preconditioning therapy | -24
fludarabine | -24
melphalan | -24
thiotepa | -24
antithymocyte globulin | -24
developed Escherichia coli sepsis | -16
started on antibiotics | -16
developed hemodynamic instability | -16
admitted to the Pediatric Intensive Care Unit | -16
developed refractory septic shock | -8
intubation | -8
volume resuscitation | -8
inotropic support | -8
venoarterial ECMO | -8
cannulated with a 14-French arterial cannula | -8
cannulated with a 14-French venous cannula | -8
echocardiogram | -8
severely diminished left ventricular function | -8
left atrial hypertension | -8
balloon atrial septostomy | -8
inotropic support weaned off | -4
required continuous renal replacement therapy | -4
received unrelated HLA donor stem cell transplant | 0
received 68 ml of ABO-mismatched cord blood transplant | 0
CD34+ count of 4.7 × 105/kg | 0
total nucleated cell count of 1.12 × 108/kg | 0
cord blood infused on the arterial side of the circuit | 0
left-sided paralysis | 72
emergent head computed tomography | 72
acute intraparenchymal hemorrhages | 72
right posterior temporal lobe | 72
left occipital lobe | 72
4 mm right to left midline shift | 72
decannulated from ECMO | 72
brain magnetic resonance | 144
stable right greater than left occipital lobe hematomas | 144
watershed infarction | 144
started to show signs of engraftment | 288
extubated | 432
fluorescence in situ hybridization XY showed 100% donor cells | 480
transitioned to peritoneal dialysis | 624
discharged to the floor | 696
discharged home | 940
peritoneal catheter removed | 954
recovered from neurologic injury | 8760
complete donor engraftment | 8760
no evidence of mixed chimerism | 8760
no signs of chronic graft versus host disease | 8760