44 years old | 0
male | 0
admitted to the hospital | 0
shortness of breath | 0
loose stools | 0
fatigue | 0
hypoxia | 0
oxygen saturations of 84% on air | 0
nonsmoker | 0
no history of previous lung disease | 0
no recent travel abroad | 0
no known contacts with SARS-CoV-2 positivity | 0
hypertension | -672
chronic glomerulonephritis | -672
stage III chronic kidney disease | -672
stable eGFR of 30–35 | -672
amlodipine | -672
doxazosin | -672
ramipril | -672
febrile | 0
dyspnoeic | 0
respiratory rate of 33/min | 0
oxygen saturation of 84% on room air | 0
septic screen | 0
intravenous antibiotics | 0
fluids | 0
urinary output monitoring | 0
patchy consolidation at the left lung base | 0
oxygen saturation of 92% on 15L of oxygen | 0
fatigue | 0
deteriorating work of breathing | 0
sedation | 0
intubation | 0
ventilation | 0
emergency transfer ventilator | 0
transferred to the ICU | 0
long term mechanical ventilation | 0
respiratory viral PCR positive for SARS-CoV-2 | 0
negative for adenovirus | 0
negative for influenza A and B | 0
negative for parainfluenza viruses | 0
negative for rhinovirus | 0
negative for human enterovirus | 0
negative urinary pneumococcal and legionella antigen testing | 0
blood-borne virus screening negative | 0
sickle cell screening negative | 0
extubated | 264
slow wean off oxygen therapy | 264
recovery | 264
physiotherapy | 264
discharged | 336
persistent exercise limiting dyspnoea | 336
malaise | 432
odynophagia | 432
anterior neck swelling | 448
persisting pain | 448
painful goitre | 448
pain on swallowing | 448
no signs of infection on examination | 448
thyrotoxicosis | 448
slight weight loss | 448
general malaise | 448
mild autonomic symptoms of heat intolerance | 448
increased resting heart rate of 90 bpm | 448
hyperthyroid picture | 448
positivity for antithyroid peroxidase antibodies | 448
raised inflammatory markers | 448
propranolol 40 mg once daily | 448
thyroid function testing | 448
ultrasound imaging of the neck | 448
geographic hypoechoic areas | 448
minimal colour flow Doppler signal | 448
reactive cervical lymph nodes | 448
normal appearance of the salivary glands | 448
no thyroid nodules | 448
hyperthyroid biochemical picture | 504
thyroid-secreting hormone 0.006 mIU/L | 504
free T4 21.7 pmol/L | 504
free T3 5.2 pmol/L | 504
anterior neck pain settled | 672
swelling and pain of the goitre reduced | 672
symptoms of thyrotoxicosis improved | 672
resolution of general malaise | 672
hot flushes | 672
corticosteroids for pain relief considered unnecessary | 672
repeat serum TSH concentration | 784
mild hypothyroid biochemical picture | 784
TSH 5.22 mIU/L | 784
hypothyroid period lasted 4 weeks | 896
normalisation of thyroid hormones | 1024