66 years old | 0
male | 0
farmer | 0
current heavy smoker | 0
96 pack-years | 0
admitted to the hospital | 0
influenza-like illness | -720
fever | -288
cough | -288
arthralgia | -288
history of pneumonia | -7200
history of acute renal failure | -14400
treated with oseltamivir | -288
high fever continued | -192
dyspnea gradually progressed | -192
admitted to a nearby hospital | -192
computed tomography scans of the chest showed bilateral multiple granular shadows and patchy opacities | -192
MRSA detected in a sputum culture | -192
treated with antibiotics | -192
C-reactive protein level reduced | -96
bilateral consolidation on chest X-ray films worsened | -96
transferred to our hospital | 0
conscious | 0
temperature 38.2 ºC | 0
blood pressure 149/79 mmHg | 0
heart rate 118 beats/minute | 0
respiratory rate 20 breaths/minute | 0
oxygen saturation 98% | 0
faint coarse crackles in the bilateral lungs | 0
no wounds observed | 0
leukocytosis with predominant neutrophils | 0
hypoalbuminemia | 0
CRP level elevated | 0
procalcitonin level 2.43 ng/mL | 0
soluble interleukin 2 receptor elevated | 0
rheumatoid factor normal | 0
antinuclear antibodies normal | 0
anticytoplasmic antibodies normal | 0
bilateral infiltration on chest X-ray film | 0
rapidly progressive formation of multiple cavities and surrounding ground-grass opacities with bilateral pleural effusion on chest CT | 0
treated with SBT/ABPC again | 0
formation of multiple cavities suggested different possible diagnoses | 0
blood culture sets negative | 0
echocardiography showed no vegetation in the cardiac valves | 0
deep vein thrombosis not observed | 0
bronchoscopy performed | 48
suctioning of purulent sputum | 48
biopsy | 48
brushing cytology | 48
gram staining showed grapelike clusters of gram-positive cocci | 48
cytological examination showed neutrophils with phagocytosis of bacterium | 48
histopathological examination showed necrosis with inflammatory exudate surrounding the neutrophils | 48
treated with VCM | 96
MRSA isolated from sputum sensitive to trimethoprim/sulfamethoxazole | 96
MRSA isolated from sputum sensitive to erythromycin | 96
MRSA isolated from sputum sensitive to minocycline | 96
MRSA isolated from sputum sensitive to clindamycin | 96
MRSA isolated from sputum sensitive to vancomycin | 96
type IV staphylococcus cassette chromosome mec identified | 96
PVL gene identified | 96
diagnosed with necrotizing pneumonia due to CA-MRSA | 96
administration of VCM reduced temperature | 96
administration of VCM reduced white blood cell count | 96
administration of VCM reduced serum level of CRP | 96
oxygenation status resolved | 96
pulmonary opacities on chest X-ray film improved | 96
changed VCM to linezolid | 648
sputum not positive for any strains of bacteria | 720
sputum not positive for MRSA | 720
discharged from the hospital | 984
chest CT scans at six months after treatment showed disappearance of multiple cavities | 4320