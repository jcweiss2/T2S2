40 years old | 0
male | 0
admitted to hospital | 0
polytrauma | -48
blunt trauma to the chest | -48
right hemothorax | -48
blunt trauma to the abdomen | -48
right lower lobe liver laceration | -48
fractured right tibia | -48
Injury severity scoring (ISS) of 26 | 0
Sequential Organ Failure Assessment (SOFA) score of 12 | 0
Acute Physiology and Chronic Health Evaluation (APACHE II) score of 18 | 0
CECT of the chest and abdomen | 0
right hemothorax | 0
right lower lobe liver laceration | 0
deranged renal parameters | 0
coagulopathy | 0
oliguric | 24
anuric | 72
sepsis | 72
multiorgan failure | 72
respiratory failure | 72
renal failure | 72
metabolic disturbance | 72
intubation | 120
ventilator support | 120
heparin-free dialysis | 72
heparin-free dialysis | 96
heparin-free dialysis | 120
no blood products transfused | 0
GCS decreased from 15 to 6 | 120
noncontrast computed tomography head | 120
massive hemorrhage in parieto-occipital region | 120
intraventricular extension | 120
surgical intervention planned | 120
coagulation profile correction planned | 120
patient expired | 126
high lactate | -48
hypovolemia | -48
contrast induced nephropathy | -48
inadequate hydration | -48
abdominal compartment syndrome | -48
myoglobinuria | -48
microvascular bleeding | 0
elevated prothrombin time (PT) | 0
elevated partial thromboplastin time (PTT) | 0
platelet dysfunction | 0
uraemia | 0
conjugated estrogens | 0
desmopressin | 0
cryoprecipitate | 0
thromboelastography (TEG) | 0