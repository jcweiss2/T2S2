39 years old | 0
    woman | 0
    diagnosed with palpable mass on her right breast | -3408
    Hodgkin lymphoma | -13632
    treated with chemotherapy | -13632
    mantle field radiation | -13632
    inflammatory colitis | -13632
    last flare | -408
    treated with mesalazine | -408
    younger sister died from metastatic myxoid liposarcoma | 0
    radiological examination of the breast | -3408
    pathological examination confirmed invasive ductal carcinoma | -3408
    triple-negative phenotype | -3408
    MIB1 85% | -3408
    staging CT scan of the thorax and abdomen | -3408
    neoadjuvant chemotherapy with paclitaxel and carboplatin | -3408
    first cycle completed | -3408
    no hematological toxicity | -3408
    port-à-cath insertion | -336
    presented to emergency room | 0
    temperature of 38.8°C | 0
    normal vital signs | 0
    subcutaneous cellulitis | 0
    colliquative necrosis | 0
    elevated white blood cell count | 0
    neutrophilia | 0
    elevated C-reactive protein | 0
    broad-spectrum i.v. antibiotic therapy | 0
    port rimotion | 0
    necrosectomy | 0
    defervescence | 0
    improvement in subcutaneous cellulitis | 0
    improvement in blood works | 0
    new febrile seizure | 96
    WBC rise | 96
    worsening of skin lesion | 96
    second necrosectomy | 96
    peripheral blood cultures negative for infection | 96
    skin plug negative for infection | 96
    i.v. catheter tip showed Klebsiella pneumoniae | 96
    antibiotic therapy modified | 96
    chest/abdomen CT scan showed mediastinitis | 96
    bilateral pleural effusion | 96
    left pulmonary atelectasis | 96
    transferred to Thoracic Surgery Unit | 96
    left thoracoscopy | 96
    pleural drainage | 96
    mediastinal drainage | 96
    admitted to Intensive Care Unit | 96
    postoperative course characterized by sepsis | 96
    required broad-spectrum antibiotic | 96
    required antifungal therapy | 96
    required hemodynamic support | 96
    required non-invasive ventilation | 96
    specimens analyzed | 96
    intensive inflammatory infiltrate | 96
    differential diagnosis included pyoderma gangrenosum | 96
    presence of triple-negative breast cancer | 96
    systemic methylprednisolone started | 96
    topical cyclosporine started | 96
    seriate chest X-ray | 96
    CT scan showed resolution of mediastinitis | 96
    resolution of pleural effusion | 96
    wound improvement with scar | 96
    normalization of blood count | 96
    normalization of flogosis index | 96
    breast ultrasound showed no change in lump dimension | 96
    multidisciplinary meeting | 96
    right mastectomy | 432
    axillary dissection | 432
    breast surgical wound healing regular | 432
    pathology assessment revealed fibroelastosis | 432
    chronic inflammation | 432
    isolated neoplastic cells | 432
    8 axillary nodes negative | 432
    restaging CT negative for distant metastasis | 432
    BRCA mutation test negative | 432
    p53 mutation test negative | 432
    released from the hospital | 528
    autologous skin graft | 528
    PICC implant | 528
    resumed chemotherapy | 528
    dose reduction | 528
    completed fourth cycle | 1344
    good tolerance | 1344
    started follow-up | 1344
    