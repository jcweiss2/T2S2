26 years old | 0
male | 0
admitted to the hospital | 0
generalized abdominal pain | -72
infrequent watery diarrhea | -72
abdominal pain radiating to flanks | -72
abdominal pain aggravating after food ingestion | -72
acute hepatitis A | -72
increased liver enzymes | -72
high HAV IgG Ab | -72
bloody diarrhea | -30
night sweats | -30
significant weight loss | -30
epigastric abdominal pain | -30
infrequent nausea/vomiting | -30
watery diarrhea | -30
stable vital signs | 0
mild epigastric tenderness | 0
splenomegaly | 0
abdominal ultrasonography | 0
moderate splenomegaly | 0
stool exam contained RBC | 0
no WBC in stool exam | 0
gastroenterologist consultation | 0
rheumatologist consultation | 0
upper gastrointestinal endoscopy | 0
chronic gastritis | 0
colon biopsy | 0
inflammatory bowel disease (IBD) | 0
fever | 24
bloody diarrhea | 24
treated by Mesalazine | 24
treated by Asacol enema | 24
treated by antibiotics | 24
peripheral blood smear (PBS) showed aggregated platelets | 48
Doppler ultrasound of the portal system | 48
portal and splenic veins with increased diameter | 48
normal flow, spectral waves | 48
normal patency of the superior mesenteric artery | 48
abdominopelvic computed tomography | 72
mesenteric fat stranding | 72
thick-walled bowels | 72
portal and superior mesenteric vein thromboses (PVT) | 72
intolerable abdominal pain | 96
generalized tenderness | 96
rebound tenderness | 96
guarding | 96
significant thrombocytopenia | 96
thrombocytopenia correction | 120
laparotomy | 120
bloody ascites | 120
colon necrosis | 120
total colectomy | 120
ileostomy | 120
mural necrosis | 120
intraluminal thrombosis of vascular canals | 120
hypotension | 144
dyspnea | 144
abnormal coagulation studies | 144
no schistocyte on PBS | 144
thrombocytopenia | 144
elevated fibrinogen | 144
elevated FDP levels | 144
treated with fresh frozen plasma | 144
death | 168
post-mortem diagnosis | 168
Factor V Leiden | 168
antiphospholipid syndrome (APS) | 168
portal system thrombosis | 168