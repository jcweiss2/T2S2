70 years old | 0
male | 0
farmer | 0
admitted to the hospital | 0
high-grade fever | -120
generalized body ache | -120
headache | -120
altered sensorium | -24
joint pains | -120
epigastric pain | -120
no comorbidities | 0
no drug addiction | 0
no intoxication | 0
inguinal lymphadenopathy | 0
mild generalized rash | 0
no eschar | 0
hemodynamically stable | 0
disoriented | 0
no focal neurological deficit | 0
no neck rigidity | 0
acute febrile illness | 0
undifferentiated fever | 0
malaria test negative | 0
dengue test negative | 0
typhoid test negative | 0
leptospira test negative | 0
scrub typhus antigen card positive | 0
scrub immunoglobulin M positive | 0
diagnosis of scrub typhus | 0
blood culture sterile | 0
body fluid culture sterile | 0
leukocytosis | 0
mild hyperbilirubinemia | 0
transaminitis | 0
slightly raised international normalized ratio | 0
hepatitis B antigen negative | 0
hepatitis C antibody negative | 0
mild fatty infiltration of the liver | 0
doxycycline treatment | 0
defervescence | 48
improved orientation | 48
weakness of lower limbs | 96
weakness progressed to upper limbs | 96
absent deep tendon reflexes | 96
flexor plantar responses | 96
bladder incontinence | 96
no bowel incontinence | 96
breathing difficulty | 96
respiratory distress | 96
intubated | 96
mechanical ventilation | 96
MRI brain normal | 96
MRI cervical spine normal | 96
nerve conduction velocity test | 96
motor sensory demyelinating polyneuropathy | 96
Guillain-Barré syndrome diagnosis | 96
cerebrospinal fluid analysis | 96
intravenous immunoglobulin therapy | 96
rifampicin treatment | 96
improvement in weakness | 168
improvement in respiratory parameters | 168
weaned off ventilator | 240
extubated | 240
oral feeding started | 240
limb physiotherapy | 240
chest physiotherapy | 240
shifted out of ICU | 240
discharged from hospital | 672
full neurological recovery | 672