67 years old | 0
Caucasian | 0
female | 0
renal transplantation | 0
deceased donor | 0
chronic renal failure | 0
unconfirmed chronic glomerulonephritis | 0
basiliximab | -672
tacrolimus | -672
mycophenolate mofetil | -672
prednisolone | -672
late onset of graft function | 0
haemodialysis dependent | 0
biopsy | -168
severe combined acute cellular rejection (2B) | -168
antibody mediated C4d positive rejection | -168
rabbit antithymocyte globulin | -168
plasmapheresis | -168
intravenous immunoglobulins | -168
recovery of graft function | -168
asymptomatic elevation of amylase | -168
asymptomatic elevation of lipase | -168
ultrasound examination (pancreas no pathology) | -168
solitary gall bladder stone | -168
conservative therapy | -168
reduced mycophenolate mofetil dose | -168
corticosteroid-dependence | -168
admitted to surgery clinic | 0
progressive sharp abdominal pain | -72
temperature > 39 C | -72
shivering | -72
tacrolimus (Advagraf) | 0
mycophenolate mofetil (Mycophenolate mofetil-SANDOZ) | 0
prednisolone (Prednison) | 0
increased serum amylase | 0
increased serum lipase | 0
normal bilirubin | 0
normal ALT | 0
normal AST | 0
normal ALP | 0
normal GGT | 0
potassium 5.3 mmol/l | 0
creatinine 384 μmol/l | 0
urea 21.9 mmol/l | 0
leukocytes 14.48 × 10^9/l | 0
CRP 433 mg/l | 0
procalcitonin 40 μg/l | 0
normal calcium | 0
normal parathyroid hormones | 0
excluded CMV | 0
excluded Epstein-Barr virus | 0
excluded herpes simplex | 0
excluded varicella zoster virus | 0
excluded acute hepatitis | 0
acute pancreatitis (CECT) | 0
subphrenic abscess collections | 0
bursa omentalis abscess | 0
fluid between small intestine loops | 0
peritonism | 0
elevated inflammatory parameters | 0
septic temperatures | 0
surgical treatment | 0
transverse laparotomy | 0
drainage of abscess subphrenically | 0
sample collection for cultivation | 0
severance of ligamentum gastrocolicum | 0
opening of bursa omentalis | 0
drainage of abscess | 0
irrigation of abdominal cavity | 0
four quadrants drainage | 0
tacrolimus discontinued | 0
mycophenolate mofetil discontinued | 0
intravenous corticoids | 0
Escherichia coli cultivation | 0
meropenem + metronidazole | 0
increased azotemia | 0
graft failure | 0
CVVHD | 0
extubation | 144
vasopressors no longer required | 144
spontaneous diuresis | 144
follow-up CECT (regression) | 216
residue after pancreas evacuation | 216
no progression of inflammatory changes | 216
regression of inflammatory parameters | 216
stabilization of laboratory values | 216
tacrolimus renewed | 72
reduced corticoids dose | 72
full sustenance | 336
surgical wound VAC system | 336
transferred to nephrological department | 336
discharged | 336
rebiopsy (no rejection) | 2160
no recurrence of acute pancreatitis | 2160
tacrolimus | 2160
prednisolone (Prednison 5 mg/day) | 2160
good graft function | 2160
