53 years old | 0
woman | 0
presented with necrotizing fasciitis | 0
transferred to ICU | 0
unconscious | 0
septic shock | 0
high temperature of 39.7°C | 0
myalgia | 0
breathing difficulties | 0
past medical history of respiratory failure | 0
past medical history of mild hypertension | 0
past medical history of obesity | 0
heavy smoker | 0
large necrotic area of skin and soft tissue | 0
purulent discharge | 0
palpable right axillary lymph nodes | 0
tachypneic | 0
heart rate of 115 bpm | 0
blood pressure of 80/50 mmHg | 0
leukocytosis | 0
increased ESR | 0
increased CRP | 0
low hemoglobin level | 0
increased serum creatine kinase | 0
resuscitated with intravenous fluids | 0
imaging performed | 0
blood samples taken | 0
treated with cefazolin | 0
treated with gentamycin | 0
hemodynamically stable | 24
underwent surgical debridement | 24
segmental partial mastectomy | 24
subtotal excision of outer quadrants of right breast | 24
nipple and areola spared | 24
intraoperative wound tissue collected | 24
exudate collected | 24
histopathological examination | 24
intubated | 24
vital signs stable | 24
hyperbaric oxygen therapy | 96
extubated | 120
Staphylococcus aureus identified | 120
Klebsiella pneumoniae identified | 120
Acinetobacter baumanii identified | 120
Staphylococcus epidermidis isolated | 120
antibiotic regimen changed to vancomycin | 120
antibiotic regimen changed to meropenem | 120
NPWT dressings applied | 24
foam dressings changed every 48 hours | 24
wounds appeared clean | 1008
pink granulation tissue present | 1008
reduced wound size | 1008
breast defect surgically repaired | 1008
nipple and areola centralization technique | 1008
defects in right chest managed with NPWT | 1008
defects in right flank managed with NPWT | 1008
discharged from hospital | 720
portable NPWT device for home use | 720
seen in clinic once a week | 720
CT scan performed every 14 days | 720
recovered well | 3360
wounds healed successfully | 3360
breast shape retained | 3360
breast volume retained | 3360
good cosmetic effect | 3360
unconscious |1 0
