29 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
admitted to hospital | 0 | 0 | Factual
muscle pain | -144 | 0 | Factual
joint pain | -144 | 0 | Factual
general weakness | -144 | 0 | Factual
fever | -144 | 0 | Factual
liver dysfunction | -144 | 0 | Factual
total bilirubin 5.7 mg/dl | -144 | 0 | Factual
serum glutamic oxaloacetic transaminase 633 U/L | -144 | 0 | Factual
serum glutamic pyruvate transaminase 412 U/L | -144 | 0 | Factual
gamma-glutamyl transferase 161 U/L | -144 | 0 | Factual
lactate dehydrogenase 1668 U/L | -144 | 0 | Factual
C-reactive protein 519 mg/l | -144 | 0 | Factual
procalcitonin 1.28 ng/ml | -144 | 0 | Factual
leukocyte levels 14.8 × 10³/μl | -144 | 0 | Factual
acute respiratory failure | 0 | 0 | Factual
altered state of consciousness | 0 | 0 | Factual
continuous sedation | 0 | 336 | Factual
muscle relaxation | 0 | 336 | Factual
intubation | 0 | 336 | Factual
mechanical ventilation | 0 | 336 | Factual
FiO2 100% | 0 | 336 | Factual
SpO2 88.7% | 0 | 336 | Factual
hemodynamic instability | 0 | 168 | Factual
norepinephrine 0.6 μg/kg/min | 0 | 168 | Factual
vasopressin not available | 0 | 0 | Factual
broad-spectrum empirical antimicrobial therapy | 0 | 168 | Factual
meropenem | 0 | 168 | Factual
azithromycin | 0 | 168 | Factual
oseltamivir | 0 | 168 | Factual
methylprednisolone | 0 | 168 | Factual
stress ulcer prophylaxis | 0 | 168 | Factual
thromboprophylaxis | 0 | 168 | Factual
CRRT | 144 | 336 | Factual
CytoSorb® | 168 | 192 | Factual
prone position | 0 | 168 | Factual
chest CT | 0 | 168 | Factual
bedside focus ultrasound | 0 | 168 | Factual
acute renal failure | 144 | 144 | Factual
septic episode | 240 | 240 | Factual
second CytoSorb® therapy | 240 | 264 | Factual
norepinephrine discontinued | 192 | 192 | Factual
inflammatory marker levels reduced | 168 | 336 | Factual
CRP decreased | 168 | 336 | Factual
leukocyte levels normalized | 168 | 336 | Factual
ICU delirium | 168 | 336 | Factual
antipsychotics | 168 | 336 | Factual
percutaneous tracheostomy | 168 | 336 | Factual
ventilator weaning | 336 | 336 | Factual
discharged from ICU | 336 | 336 | Factual
transferred to general ward | 336 | 336 | Factual
transferred to rehabilitation clinic | 360 | 360 | Factual
influenza A (H1N1) | -144 | 0 | Factual
bilateral pneumonia | -144 | 0 | Factual
massive bilateral pneumonia | 0 | 168 | Factual
minimal pleural effusions | 0 | 168 | Factual
lung-protective ventilation | 0 | 336 | Factual
control of inflammatory response | 168 | 336 | Factual
hemodynamic stabilization | 168 | 336 | Factual
decrease in inflammation markers | 168 | 336 | Factual
improvement in patient ventilation parameters | 168 | 336 | Factual
improvement in lung function | 168 | 336 | Factual
decrease in vasopressors | 168 | 336 | Factual