46 years old | 0  
    male | 0  
    referred to the hospital | 0  
    sudden pain | 0  
    redness | 0  
    hardening in the lateral side of the left thigh | 0  
    subfebrile fever | 0  
    no anamnesis of trauma/injury | 0  
    no immunosuppression | 0  
    right thigh pain | -2160  
    recurrent episodes of lateral side of left thigh pain | -336  
    swelling | -336  
    worsened in the last 24 hours | -24  
    relapsed to pneumonia | -4320  
    onset of the first symptoms of osteomyelitis | -4320  
    no evidence of immunosuppression | 0  
    mild leukocytosis | 0  
    significant thrombocytosis | 0  
    moderately elevated C-reactive protein | 0  
    normal blood biochemistries | 0  
    normal urine analysis | 0  
    increased partial CO2 | 0  
    X-ray showing left femoral destruction | 0  
    CT scan showing abscess in the left thigh | 0  
    symptoms recurred | 2160  
    pathologic fracture of the left femoral diaphysis | 2160  
    displacement | 2160  
    osteomyelitis of the left femur | 2160  
    osteomyelitis of the right femur | 2160  
    sequester | 2160  
    contrast flow around the implant | 2160  
    air inserts in interfascial spaces | 2160  
    abscess in the intramedullary space in the right femur | 2160  
    fistulas merging with the intramedullary space | 2160  
    bone destruction | 2160  
    abscess around the femur | 2160  
    destructive processes in the left femur | 2160  
    longitudinal air inserts in the interfascial space | 2160  
    pathological fracture in the right femur | 4320  
    right femur completely healed | 8640  
    external AO fixation | 2160  
    left femur shortening by 5 cm | 8640  
    Anaerococcus prevotii identified | 0  
    sensitive to ampicillin and penicillin | 0  
    lung infiltrates | 0  
    purulent processes on the molars | 0  
    mixed microflora | 0  
    spontaneous reciprocal haematogenous osteomyelitis of the femurs | 0  
    secondary abscesses on both thighs | 0  
    sepsis | 0  
    abscessotomy | 0  
    active wash | 0  
    antibiotics treatment | 0  
    debridement surgery | 0  
    postoperative wound excision | 2160  
    femoral trepanation | 2160  
    regular washes | 2160  
    external osteosynthesis of the left femur | 2160  
    preventive external AO fixation on the right femur | 2160  
    pathological fracture without displacement of the right femur | 4320  
    AO switched to external fixation with Ilizarov's apparatus | 4320  
    condition worsened | 8640  
    secretion around the bars | 8640  
    severe pain of the left thigh | 8640  
    re-inoculation | 8640  
    treatment with intramedullary necklace of antibiotics | 8640  
    external fixation with Ilizarov's apparatus again | 8640  
    condition improved | 12960  
    removal of the proximal ring on the left side | 12960  
    redness of the left thigh | 17520  
    intense pain | 17520  
    febrile fever | 17520  
    purulent discharge around the bars | 17520  
    four operations | 17520  
    debridements | 17520  
    intramedullary osteosynthesis with silver-plated nail | 17520  
    long-term antibiotic therapy with Meropenem and Penicillin | 17520  
    left knee remodeling | 17520  
    passive knee motion machine | 17520  
    left leg radiographically shorter by 5 cm | 17520  
    intense left knee and thigh pain | 21840  
    protrusion of a protruding propellant through the skin | 21840  
    extensive wound secretion | 21840  
    migration of the screws | 21840  
    screw pierced the skin | 21840  
    operative treatment - abscessotomy | 21840  
    crop | 21840  
    biopsy | 21840  
    pathological examination | 21840  
    instability of the intramedullary nail | 21840  
    distal femur fixed by external fixation | 21840  
    removal of the intramedullary nail | 21840  
    removal of external fixation apparatus | 21840  
    debridement on the left thigh | 21840  
    repeated debridement | 24000  
    constant washing | 24000  
    no improvement | 24000  
    debridement | 24000  
    external fixation with Ilizarov's apparatus | 24000  
    four reconstructive/plastic surgeries of the left thigh | 24000  
    transplantation of free fibula into femur | 24000  
    postoperative period complicated by infectious complication | 24000  
    purulent secretion from the wound | 24000  
    fistula | 24000  
    amputation of the left femur | 24000  
    sepsis complication | 24000  
    treatment in the intensive care unit | 24000  
    stump debridement | 24000  
    Meropenem | 24000  
    Colistin | 24000  
    right femur healed completely | 28800  
    signs of osteomyelitis did not appear | 28800  
    positive clinical effects on the stump | 28800  
    stump healed | 28800  
    discharged in satisfactory condition | 28800  
    rehabilitation treatment | 28800  
    outpatient follow-up for about a year | 28800  
    all signs of osteomyelitis disappeared | 28800  
