60 years old|0
male|0
alcohol abuse|0
hypertension|0
hydrochlorothiazide|0
admitted to the hospital|0
acute delirium|0
Methicillin-sensitive Staphylococcus aureus (MSSA) bacteremia|0
aortic valvular endocarditis|0
disseminated septic emboli|0
MSSA meningitis|0
C6-7 osteomyelitis|0
spinal abscess|0
sternoclavicular joint abscess|0
multiple septic emboli infarcts in the brain|0
multiple septic emboli infarcts in the liver|0
multiple septic emboli infarcts in the spleen|0
multiple septic emboli infarcts in the kidneys|0
aortic valve replacement|0
significant upper gastrointestinal (GI) bleeding|0
aggressive blood transfusions|0
duodenal ulcers with visible vessels|0
endoscopy|0
active bleeding on five subsequent endoscopies|0
epinephrine injection|0
BICAP cauterization|0
endoclipping of vessels|0
hemospray with procoagulant|0
argon plasma coagulation|0
IR embolization of the gastroduodenal artery|0
IR embolization of multiple branches of the superior pancreaticoduodenal arteries|0
IR embolization of multiple branches of the inferior pancreaticoduodenal arteries|0
continued hemorrhage|0
daily transfusions|0
hemodynamic stability|0
generalized mucosal bleed throughout the duodenum|0
duodenal resection|0
Whipple procedure|0
unrelenting duodenal hemorrhage|0
high risk for pancreaticojejunostomy anastomotic leak|0
high mortality risk|0
duodenal resection with total pancreatectomy|0
duodenal resection with splenectomy|0
multiple aberrant blood vessels extending into the duodenum|0
critically ill|0
transfer to ICU|0
gastrojejunostomy|24
hepaticojejunostomy|24
flattened duodenal mucosa|0
congested duodenal mucosa|0
focally ulcerated duodenal mucosa|0
viral cytopathic changes|0
autolysis of duodenal mucosa|0
no vasculitis|0
no intravascular thrombi|0
patchy panlobular coagulative necrosis in pancreas|0
non-occlusive thrombi within muscularized arteries|0
viral cytopathic changes in ductal epithelial cells|0
immunohistochemical stains for CMV positive in duodenum|0
immunohistochemical stains for CMV positive in pancreas|0
mild reactive gastropathy|0
no Helicobacter gastritis|0
nonreactive CMV IgM antibodies|0
reactive CMV IgG antibodies|0
negative DNA quantitative PCR for CMV|0
normal HIV immunologic assays|0
normal hepatitis B immunologic assays|0
normal hepatitis C immunologic assays|0
hemodynamically stable|72
no additional blood transfusions|72
intravenous ganciclovir|72
oral valganciclovir|168
monitoring for pancytopenia|168
monitoring for renal dysfunction|168
monitoring for CMV reactivation|168
no history of immunosuppressive treatments|0
no history of immunosuppressive infections|0
transient depression in immunity|0
ICU admission|0
use of antibiotics|0
use of antacids|0
use of H2 blockers|0
use of PPIs|0
risk factors for CMV reactivation|0
severe necrotizing acute pancreatitis|0
autolysis of duodenal mucosa by pancreatic juice|0
