48 years old | 0
female | 0
admitted to the emergency department | 0
complaining of left breast enlargement | 0
black discoloration of breast skin | 0
fever | -8760
loss of appetite | -8760
weight loss | -8760
diabetes mellitus | -8760
hypertension | -8760
no previous history of lymphoma | 0
no previous history of breast implant | 0
no family history of breast cancer | 0
no family history of lymphoma | 0
left breast swollen | 0
dark discoloration of breast skin | 0
multiple small punched-out ulcers | 0
discharging purulent material | 0
nipple retracted | 0
breast tender | 0
breast warm | 0
breast firm | 0
large palpable left axillary lymph node | 0
marked leukocytosis | 0
prolongation of coagulation profile markers | 0
microbiological cultures positive for MRSA | 0
emergency surgery | 0
simple mastectomy | 0
died 2 days after operation | 48
disseminated intravascular coagulation | 48
septicemia secondary to MRSA | 48
no autopsy study | 48
mastectomy specimen received | 0
black ulcerated gangrenous skin | 0
retracted nipple | 0
multiple firm tan-white focally necrotic solid tumor nodules | 0
tumor cells with ample eosinophilic to amphophilic cytoplasm | 0
nuclear pleomorphism | 0
coarsely clumped chromatin pattern | 0
irregular nuclear membrane | 0
basophilic micro- and macronucleoli | 0
hallmark cells | 0
wreath-like appearance | 0
bizarre nuclear shapes | 0
mummified cells | 0
Reed-Sternberg cells-like morphology | 0
emperipolesis | 0
brisk mitotic activity | 0
atypical mitotic figures | 0
mixed inflammatory cell infiltrate | 0
perivascular distribution of tumor cells | 0
un-involved atrophic ducts and lobules | 0
focal ulcerations | 0
no epidermotropism | 0
perineural invasion | 0
tumor cells positive for CD30 | 0
tumor cells positive for CD45 | 0
tumor cells positive for CD45RO | 0
tumor cells positive for granzyme B | 0
tumor cells positive for TIA-1 | 0
tumor cells positive for vimentin | 0
tumor cells positive for CD4 | 0
tumor cells positive for CD43 | 0
tumor cells positive for EMA | 0
tumor cells positive for BCL-6 | 0
tumor cells positive for BCL-2 | 0
loss of CD1a | 0
loss of CD3 | 0
loss of CD5 | 0
loss of CD8 | 0
loss of CD7 | 0
loss of CD2 | 0
loss of CD20 | 0
loss of CD19 | 0
loss of CD79a | 0
loss of PAX-5 | 0
loss of ALK-1 | 0
loss of CD15 | 0
loss of CD68 | 0
loss of pancytokeratins | 0
loss of S100 protein | 0
loss of desmin | 0
loss of SMA | 0
loss of HMB-45 | 0
loss of P63 | 0
loss of E-cadherin | 0
high MIB-1 labeling index | 0
diagnosis of PB-ALCL, giant cell-rich pattern | 0