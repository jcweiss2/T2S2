48 years old | 0
    woman | 0
    long-standing history of intractable migraine headaches | 0
    admitted to specialty headache unit | 0
    aggressive management | 0
    no known history of peripheral vascular disease | 0
    no known history of cardiac disease | 0
    multiple admissions for treatment of headaches since 2003 | 0
    received dihydroergotamine mesylate (DHE) 45 during previous hospitalizations | 0
    received two courses of DHE 0.5 mg × 1 | 0
    received 1 mg every 8 h for total of eight doses on days 1–3 | 0
    second course of therapy on days 7–9 | 0
    became obtunded | 96
    became minimally responsive | 96
    became hypotensive | 96
    blood pressure 80/45 mm Hg | 96
    abdomen moderately distended | 96
    few bowel sounds | 96
    lactate acid level 4.5 mmol/l | 96
    white blood cell count 18.0 | 96
    17% bands | 96
    stool Clostridium difficile negative | 96
    transferred to intensive care unit | 96
    given intravenous fluid boluses | 96
    started on vasopressors | 96
    given broad spectrum antibiotics | 96
    eventually required intubation | 96
    chest radiograph unremarkable | 96
    abdominal x-rays showed mild prominence of the colon | 96
    became progressively acidotic | 96
    worsening bandemia | 96
    colonoscopy showed diffuse ischemic colitis | 96
    fecal impaction | 96
    no pseudomembranes | 96
    taken to operating room | 96
    underwent laparotomy | 96
    peritoneal cavity filled with murky, foul-smelling fluid | 96
    gangrene of the descending colon | 96
    necrosis distal to splenic flexure to sigmoid colon | 96
    large amount of impacted stool in left colon | 96
    vasculature intact with audible Doppler signals | 96
    removal of gangrenous bowel | 96
    condition improved promptly | 96
    final pathology showed 86 cm of patchy, dark green/black large bowel | 96
    consistent with ischemic necrosis | 96
    bowel wall intact throughout | 96
    final diagnosis of gangrenous large bowel | 96
    ischemic colitis | 96
    thrombi or emboli noted | 96
    hypercoagulable panel performed | 96
    negative for clotting disorders | 96
    no history of cardiac arrhythmias | 0
    non-smoker | 0
    no cardiac risk factors | 0
    no history of post-prandial pain | 0
    no food fear | 0
    no signs of venous congestion | 96
    no signs of stasis at surgery | 96
    no hypercoagulable disorder | 96
    colon not edematous | 96
    no clot identified in vasculature | 96
    most probable cause: non-occlusive mesenteric ischemia | 96
    left colic artery vasoconstriction induced by ergotamine | 96
    bowel wall distention from impacted stool | 96
    DHE dosing exceeding recommendations | 0
    received 17 mg DHE over 9 days | 0
    ischemic colitis secondary to high-dose ergotamine | 96
    fourth reported case of ischemic colitis secondary to ergotamine | 96
    first requiring colon resection | 96
    patient informed of risks of ischemia | 96
    ischemic colitis considered in differential diagnosis | 96
    