33 years old| 0
    woman| 0
    childhood history of hydronephrosis| 0
    hydronephrosis secondary to vesicoureteral reflux| 0
    vesicoureteral reflux| 0
    9-year history of erythroderma| -94896
    confluent folliculocentric erythematous scaly plaques| -94896
    islands of sparing| -94896
    orange palmoplantar hyperkeratosis| -94896
    eczematous lesions| -94896
    differential diagnoses| 0
    PRP| 0
    psoriasis| 0
    atopic dermatitis| 0
    epidermotropic cutaneous T-cell lymphoma| 0
    search for skin and blood T-cell clone| 0
    negative T-cell clone| 0
    blood screening| 0
    no Sezary cells| 0
    no phenotypically atypical lymphocytes| 0
    whole genome sequencing| 0
    CARD14 sequencing| 0
    no causal mutation found| 0
    skin biopsy specimens| 0
    epidermal acanthosis| 0
    alternating orthokeratosis and parakeratosis| 0
    dermal lymphohistiocytic infiltrate| 0
    few neutrophils| 0
    type II PRP diagnosed| 0
    severe clinical course| 0
    intense erythroderma| 0
    Staphylococcus aureus septicemia| 0
    two admissions in intensive care unit| 0
    severe depression| 0
    anorexia| 0
    loss of 30 kg| 0
    previous unsuccessful treatments| -8784
    topical corticosteroids| -8784
    acitretin| -8784
    photochemotherapy| -8784
    cyclosporine| -8784
    methotrexate| -8784
    infliximab| -8784
    ustekinumab| -8784
    intravenous immunoglobulin| -8784
    omalizumab| -8784
    prednisone efficient| -8784
    relapse with less than 0.5 mg/kg/d prednisone| -8784
    condition partially improved with cyclosporine (5 mg/kg/d)| 0
    cyclosporine association| 0
    10 mg prednisone| 0
    informed consent| 0
    secukinumab initiated| 0
    association with cyclosporine| 0
    association with 10 mg prednisone| 0
    received 5 subcutaneous 300-mg weekly injections| 0
    once-a-month injections| 168
    significant clinical response after 4 weeks| 672
    prompt clinical response| 672
    quality-of-life improvement| 672
    psoriasis area and severity index decreased| 672
    dermatologic life quality index score decreased| 672
    secukinumab well tolerated| 672
    oral and esophageal candidiasis| 672
    treated with fluconazole for 14 days| 672
    secukinumab effective on clinical symptoms| 672
    quality of life improvement| 672
    no recurrence of PRP lesions with 6-month follow-up| 4320
    pruritus relief after 1 week of treatment| 168
    improvement of erythematous plaques after 2 weeks of treatment| 336
    improvement of palmoplantar keratoderma after 2 weeks of treatment| 336
    