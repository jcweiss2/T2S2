51 years old | 0
male | 0
motorcycle accident | -1
hemodynamic instability | 0
pelvic fracture | 0
soft tissue injury | 0
scrotum injury | 0
perineum injury | 0
anus injury | 0
absence of anal reflex | 0
extended EcoFast | 0
no fluid collection in abdomen | 0
no pneumothorax | 0
pelvis X-ray | 0
ischiopubic fracture | 0
ileopubic fracture | 0
symphyseal disruption | 0
resuscitation phase | 0
full-body computed tomography (CT) | 1
transfer to operating theater | 1
external screws | 2
exploratory laparotomy | 2
loop colostomy | 2
admitted to ICU | 2
no bowel function | 2
abdominal distension | 166
elevated inflammatory indices | 166
fever | 166
abdominal CT | 166
intestinal obstruction | 166
dilated small bowel loops | 166
air/fluid levels | 166
ileum segment trapped in sacral fracture | 166
exploratory laparotomy | 170
small bowel resection | 170
end-to-end manual anastomosis | 170
discharged from ICU | 200
evaluation of rectal sphincter | 200
normal rectal sphincter function | 200
colostomy closure | 210
peroneal wound healed | 210