79 years old | 0
female | 0
admitted to the hospital | 0
dyspnea | 0
palpitations | 0
no chest pain | 0
hypertension | -8760
type 2 diabetes mellitus | -8760
atrial fibrillation | -8760
colonic diverticulosis | -8760
depressive syndrome | -8760
osteoporosis | -8760
mastectomy | -2628
breast cancer | -2628
ischemic cardiomyopathy | -1752
acute myocardial infarction | -1752
percutaneous angioplasty | -1752
omeprazole | -720
metformin | -720
calcifediol | -720
calcium | -720
alendronate | -720
acenocumarol | -720
amiodarone | -720
torasemide | -720
enalapril | -720
letrozole | -720
citalopram | -720
acetaminophen | -720
lormetazepam | -720
pale | 0
diaphoretic | 0
hypothermic | 0
tachycardia | 0
aortic murmur | 0
chronic venous insufficiency | 0
no edemas | 0
hypophonesis | 0
crackles | 0
cardiac insufficiency | 2
atrial fibrillation | 2
fast ventricular response | 2
diuretics | 2
vasodilators | 2
digoxin | 2
apical and mid-segment akinesia | 2
hypokinesis | 2
myocardial damage | 2
elevated cardiac troponin | 2
leucocytosis | 2
increased inflammatory markers | 2
vascular redistribution | 2
cardiomegaly | 2
pulmonary edema | 2
coronary angiography | 2
no stenotic changes | 2
ventriculography | 2
apical dyskinesia | 2
Takotsubian apical ballooning | 2
preserved LVEF | 2
transdermal nitrates | 2
decrease in myocardial damage markers | 120
electrocardiographic stability | 120
normofrequent atrial fibrillation | 120
hyperthyroidism | 120
thyrotropin | 120
free thyroxine | 120
no goiter | 120
no exophthalmos | 120
no pretibial myxedema | 120
antibody study | 120
thyroid-stimulating immunoglobulin | 120
anti-thyroperoxidase | 120
anti-thyroglobulin | 120
amiodarone-induced hyperthyroidism | 120
methimazole | 120
ineffective treatment | 144
prednisone | 144
good response | 168
thyrotropin | 168
free thyroxine | 168
free triiodothyronine | 168
ischemic colitis | 168
bowel perforation | 168
right hemicolectomy | 168
corticoids | 168
normal thyroid function | 432
complete resolution of TC | 432
cardiovascular symptoms | 432
baseline situation | 432
new episode of ischemic colitis | 2160
bowel perforation | 2160
generalized sepsis | 2160
fatal outcome | 2160
normal thyroid function | 2160