28 years old | 0
woman | 0
8 weeks pregnant | 0
acute severe asthma | 0
short non-infective prodrome | 0
hypoxic cardiac arrest | 0
ventricular fibrillation | 0
resuscitation | 0
sinus tachycardia | 0
endotracheal intubation | 0
transfer to ICU | 0
therapeutic cooling to 33°C | 0
salbutamol (inhaled) | 0
salbutamol (intravenous) | 0
ipratropium | 0
aminophylline | 0
hydrocortisone | 0
magnesium | 0
ketamine | 0
inhalation anesthesia with 1 MAC isoflurane | 0
severe hypercapnic acidosis | 0
inadequate minute ventilation | 0
neuromuscular blockade | 0
ventilation improving | 48
ceased intravenous sedatives | 48
ceased neuromuscular blockade | 48
0.25–0.5 MAC isoflurane | 48
generalised status myoclonus | 48
stopped isoflurane | 96
comatose | 96
absent motor response to painful stimulus | 96
preserved pupillary reflexes | 96
preserved corneal reflexes | 96
preserved cough reflexes | 96
preserved gag reflexes | 96
spontaneously breathing | 96
severe generalised status myoclonus | 96
refractory to three antiepileptic medications | 96
generalised periodic discharges | 96
no discernable background rhythm | 96
reversible causes of coma eliminated | 96
clinical examination | 96
specific investigations | 96
duration of action of sedative medications | 96
no agreement about neurological outcome | 192
interethnic marriage | 192
pregnancy | 192
intensive social work support | 192
delayed onset of GSM at 48 h | 192
plasma neuron-specific enolase 51 mcg/L | 240
somatosensory-evoked potential unhelpful | 240
brain MRI performed | 240
bilateral basal ganglia infarction | 240
frontoparietal cortex infarction | 240
medical consensus regarding poor prognosis | 240
extubated | 240
died | 264
