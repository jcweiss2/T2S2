70 years old | 0
male | 0
hypertension | 0
diabetes |&nbsp;0
auricular fibrillation | 0
adenocarcinoma of the sigmoid colon stage T4aN1M0 | 0
laparoscopic exploration | 0
perforated neoplasm of the sigma infiltrating terminal ileum and right colon | 0
open surgery | 0
total oncologic colectomy | 0
ileo-rectal stapled anastomosis | 0
self-limited abdominal bleeding | 48
high dose of low molecular weight heparin | 48
hiccups | 48
haloperidol | 48
chlorpromazine | 48
CT scan | 48
absence of intraabdominal complication | 48
admitted to intensive care unit | 48
fever peaks | 72
bacteraemia related to CVC | 72
inflammatory signs on the right jugular venous access | 72
cervicothoracic CT | 72
thrombus | 72
air bubbles into the right jugular vein | 72
dilatation of an area of the vein intimately related to the phrenic nerve | 72
persistent hiccups secondary to septic thrombosis of the jugular vein | 72
treatment with LMWH | 72
antibiotics | 72
catheter removal raised doubts | 72
discharged from intensive care unit to surgery ward | 168
isolated fever peaks | 192
catheter removal | 192
3 weeks’ intravenous antibiotic cycle | 504
discharged from the hospital | 504
