28 years old | 0
male | 0
homeless | 0
Nepalese | 0
immigrated to the United States | -6*24
productive cough | -432
weight loss | -432
intermittent abdominal pain | -432
admitted to the hospital | 0
grade 3/6 systolic murmur | 0
elevated hepatic transaminases | 0
bilateral pleural effusions | 0
normal abdomen and pelvis CT | 0
general surgery consultation | 0
infectious disease consultation | 0
no antibiotics | 0
no surgical intervention | 0
transthoracic echocardiogram | 0
normal ejection fraction | 0
mobile vegetation attached to the pulmonary valve | 0
pulmonary insufficiency | 0
elevated right heart pressures | 0
bulky lesions attached to the aortic valve | 0
moderate to severe aortic insufficiency | 0
cardiogenic shock | 168
septic shock | 168
acute hypoxic respiratory failure | 168
treated with intravenous vancomycin | 168
treated with ceftriaxone | 168
transferred to a tertiary care facility | 168
multi-organ failure | 168
increased serum lactate level | 168
worsening oliguria | 168
initiation of continuous renal replacement therapy | 168
medically stabilize the patient | 168
serology testing | 0
molecular testing | 0
QuantiFERON-TB Gold In-Tube testing | 0
latent tuberculosis infection | 0
chest x-ray findings not consistent with active pulmonary tuberculosis | 0
three sputum specimens negative for acid-fast bacilli | 0
Bartonella henselae IgM positive | 0
Bartonella henselae IgG positive | 0
Bartonella quintana IgM positive | 0
Bartonella quintana IgG positive | 0
intravenous doxycycline treatment | 312
intravenous gentamicin treatment | 312
Candida albicans grown | 1440
treated with intravenous micafungin | 1440
mechanical aortic valve replacement | 1032
mitral valve repair | 1032
16S ribosomal RNA polymerase chain reaction testing | 1032
positive for Bartonella quintana | 1032
histopathology of the aortic valve | 1032
histopathology of the pulmonary valve | 1032
vegetations and destruction of the valve tissue | 1032
fibrinoid necrosis and inflammation | 1032
Warthin-Starry silver stain negative | 1032
peri-aortic thrombosis | 1200
surgical wound dehiscence | 1200
multiple thoracotomies | 1200
postoperative hemothorax | 1440
gastrointestinal bleeding | 1440
hemorrhagic shock | 1440
died | 1440