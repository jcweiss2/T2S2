62 years old | 0
female | 0
end-stage renal disease | -5760
haemodialysis | -5760
double-lumen tunnelled catheter | -5760
shortness of breath | -72
cough | -72
admitted to the emergency department | 0
tachypneic | 0
temperature 37.7° C | 0
heart rate 110 beats per minute | 0
blood pressure 100/55 mm Hg | 0
oxygen saturation 85% | 0
pansystolic murmur | 0
CT pulmonary angiography | 0
bilateral segmental and subsegmental pulmonary embolism | 0
intravenous heparin infusion | 0
hypotension | 48
ST-segment elevation | 48
elevated cardiac enzymes | 48
dilated right side | 48
significant tricuspid regurgitation | 48
normal aortic valve | 48
coronary angiography | 48
total occlusion of the posterior descending artery | 48
complete heart block | 96
temporary pacemaker insertion | 96
feverish | 96
pus oozing from the haemodialysis catheter site | 96
line sepsis | 96
catheter removal | 96
Methicillin-resistant Staphylococcus aureus | 96
transesophageal echocardiography | 96
aortic valve vegetations | 96
acute severe aortic regurgitation | 96
right atrial appendage mass | 96
patent foramen ovale | 96
intravenous vancomycin | 96
disturbed level of consciousness | 102
resistant shock | 102
mechanical ventilation | 102
intravenous inotropes | 102
extracorporeal membrane oxygenation | 102
death | 102