42 years old | 0
male | 0
admitted to the hospital | 0
severe bilateral lower extremity pain | -504
constant bilateral lower extremity pain | -504
bilateral lower extremity pain located at upper thighs | -504
radiation down the legs | -504
non-radiating severe frontal throbbing headache | -168
headache associated with occasional episodes of diplopia | -168
no stiff neck | 0
no photophobia | 0
bilateral lower extremity weakness | -96
inability to walk | -96
inability to stand | -96
nausea | 0
vomiting | 0
low-grade fever of 37.7°C | 0
no recent travel abroad | 0
no sick contacts | 0
no medical problems | 0
no previous surgical interventions | 0
20 pack year history of smoking | 0
chronic alcohol intake of four 8 oz cans of beer daily for twenty years | 0
construction worker | 0
vital signs stable on admission | 0
somnolent but arousable | 0
no acute distress | 0
unremarkable neurological examination | 0
hypereflexia of right brachioradialis | 0
hypereflexia of right biceps | 0
decrease of muscle strength in bilateral lower extremities | 0
unremarkable physical examination of other body systems | 0
mild hyponatremia | 0
mild transaminase elevation | 0
hyperbilirubinemia | 0
ammonia level in upper normal range | 0
negative urinalysis | 0
negative urine toxicology screen | 0
negative alcohol level | 0
negative hepatitis serology panel | 0
negative HIV | 0
unremarkable chest x-ray | 0
CT brain revealing multiple intraaxial hyperdense lesions with surrounding vasogenic edema | 0
chest-CT demonstrating bilateral cavitary nodules | 0
chest-CT demonstrating right hilar lymphadenopathy | 0
empiric antibiotics started: vancomycin | 0
empiric antibiotics started: ceftriaxone | 0
dexamethasone for cerebral edema | 0
MRI brain revealing multiple bilateral rim enhancing lesions | 24
negative blood cultures | 0
negative urine cultures | 0
pulmonary service consulted for bronchoscopy | 24
bronchoscopy revealing normal airway anatomy | 24
diffusely erythematous mucosa | 24
clear secretions | 24
BAL obtained from left upper lobe | 24
BAL cytology report no significant findings | 24
BAL cultures negative for fungal | 24
BAL cultures negative for bacteria | 24
BAL cultures negative for mycobacteria | 24
AFB stain negative | 24
infectious disease service consulted | 24
PPD test negative | 24
QuantiFERON Gold negative | 24
coccidioid serology negative | 24
aspergillus antigen negative | 24
toxoplasma IgG antibody negative | 24
serum cryptococcal antigen negative | 24
lumbar puncture performed | 24
CSF analysis elevated WBC count | 24
CSF appearance clear and colorless | 24
CSF neutrophils 64% | 24
CSF lymphocytes 25% | 24
CSF monocytes 11% | 24
CSF protein 37 mg/dL | 24
CSF glucose 55 mg/dL | 24
CSF serology negative | 24
CSF culture negative | 24
echocardiogram no vegetations | 24
neurosurgery consulted for brain biopsy | 24
brain biopsy not possible | 24
mental status deteriorated to disoriented to time and place | 240
oriented to person | 240
weakness of left upper extremity | 288
unsteady antalgic gait | 288
right upper extremity weakness | 312
ptosis | 312
right lower facial weakness | 312
cardiothoracic surgery consulted for VATS biopsy | 312
lung lesion unsuitable for surgical access | 312
GCS decreased to 7 | 360
bradycardic | 360
complete right sided paralysis | 360
positive right side Babinski | 360
transferred to MICU | 360
repeat head-CT with contrast revealing multiple ring enhancing lesions | 360
amphotericin B started | 360
antibiotics continued | 360
dexamethasone continued | 360
tachycardic (HR 120@130 bpm) | 456
desaturation <80% | 456
intubated | 456
mechanical ventilation support | 456
albendazole started | 456
pyrimethamine started | 456
sulfadiazine started | 456
leucovorin started | 456
continued fevers 38.7°C to 39°C | 456
clinical status worsening | 456
tissue biopsy attempts continued | 456
patient expired on twentieth hospital day | 480
autopsy performed | 528
bilateral serosanguineous pleural effusions | 528
lung abscess at right hilum | 528
microabscess formation in right hilum abscess | 528
multiple bilateral cavities in brain | 528
Gram positive branching rods in abscesses | 528
nocardia species cultured | 528
PCR analysis revealing nocardia wallacei | 528
resistance to ceftriaxone | 528
resistance to levofloxacin | 528
resistance to aminoglycosides | 528
resistance to sulfonamides | 528
sensitivity to imipenem | 528
final autopsy diagnosis nocardia pneumonitis and encephalitis | 528
cause of death systemic nocardiosis | 528
