57 years old | 0
mechanic | 0
medical history of occasional use of cocaine | 0
gradually worsening vision | -29280
optic nerve atrophy | -29280
tripped over a low brick wall | -29280
fell about one meter on the back of his head | -29280
tetraplegic | 0
transferred to a level 1 trauma center | 0
complete cord lesion on the level of C3 and C4 | 0
computed tomography showed congenital narrowing of the spinal canal at the level of C3 and C4 | 0
old fracture of the third thoracic vertebra | 0
magnetic resonance scanning showed hemorrhage in the myelum at the level of C3 and C4 | 0
transferred to the Intensive Care Unit | 0
ventilator support | 0
acute respiratory distress syndrome (ARDS) | 72
pneumonia in the right lower lobe | 72
aspiration | 72
purulent sputum removed repeatedly | 72
sputum grew Haemolytic Streptococcus group C | 72
sputum grew Streptococcus pneumoniae | 72
sputum grew Haemophilus influenzae | 72
sputum grew Enterobacter cloacae | 72
treated with piperacillin/tazobactam | 72
percutaneous tracheostomy | 240
weaning was possible | 240
no longer dependent on ventilator support | 480
spent 32 days on the Intensive Care Unit | 768
discharged to a rehabilitation center | 76 days (not converted to hours as time is already relative)
admitted again to the department of Internal Medicine | 1824
fever | 1824
diarrhea | 1824
productive cough | 1824
radiology suspect for pulmonary tuberculosis | 1824
Mycobacterium tuberculosis found in gastric contents | 1824
placed on tuberculostatic triple therapy | 1824
pseudomembranous colitis caused by Clostridium toxins | 1824
given metronidazol | 1824
free of diarrhea after ten days | 1824+240=2064
deep venous thrombosis in the right subclavian vein | 2064
erysipelas | 2064
ulceration on the fingers | 2064
cultured Escherichia coli | 2064
cultured Klebsiella pneumoniae | 2064
cultured Pseudomonas aeruginosa | 2064
cultured Morganella morganii | 2064
cultured Proteus mirabilis | 2064
urine positive for Klebsiella pneumoniae | 2064
urine positive for Enterococcus faecalis | 2064
ulcers treated surgically | 2064
heterozygosity in MBL2 exon 1 (AC genotype) | 0
heterozygosity in MBL2 promoter region Y-221X (YX genotype) | 0
homozygosity for the minor allele in MASP2 Y371D (DD genotype) | 0
heterozygosity in FCN2 T236M (TM genotype) | 0
heterozygosity in FCN2 A258S (AS genotype) | 0
homozygosity for the minor allele in TLR2 T-16934A (AA genotype) | 0
heterozygosity in CD14 C-159T (CD genotype) | 0
magnetic resonance scanning showed hemorrhage in the myelum at the level of C3 and C4 |@0
