40 years old | 0
Asian | 0
male | 0
parotid cancer | -8760
metastatic to brain | -8760
metastatic to lung | -8760
metastatic to liver | -8760
metastatic to bone | -8760
radiation | -8760
chemotherapy | -8760
palliative whole brain radiation | -8760
urinary retention | 0
ascending paralysis | 0
MRI | 0
spinal tumor | 0
emergent XRT to spine | 0
upper body weakness | 3
respiratory distress | 3
intubation | 6
cognitively intact | 6
wife arrived | 24
discussed prognosis | 24
elective intubation | 24
stated "I want to die today" | 48
restated wishes | 48
wife requested privacy | 48
changed mind | 72
wanted to live as long as possible | 72
feeding tube | 96
tracheotomy | 96
postoperative course complicated | 96
pneumonia | 120
hypotension | 120
sepsis | 120
intensive care | 120
stated "I want to die" again | 456
advocated to honor wishes | 456
wife believed patient was confused | 456
patient stated "I want you to take away the tube and let me die" | 504
family meeting | 504
wife did not agree to extubation | 504
patient's condition deteriorated | 576
became confused and agitated | 576
wife requested withdrawal of life support | 576
transferred to private room | 576
extubation | 576
died peacefully | 578