73 years old | 0
female | 0
admitted to the hospital | 0
axial diaphragma hernia | -8760
sigma diverticulosis | -8760
atrial flutter | -24
fatigue | -24
dizziness | -24
dyspnoea | -24
rapid regular pulse rate | -24
normal lung and heart sounds | -24
no peripheral oedema | -24
unclear mass on the anterior right atrial wall | -24
heterogeneous, isoechoic, immobile mass | -24
circular, hypoechoic pericardial effusion | -24
compression of the right atrium | -24
pericardiocentesis | -24
tumour screening | -24
computed tomography of skull, abdomen, thorax, and pelvis | -24
endoscopy of the upper and lower gastrointestinal tract | -24
dermatologic and gynaecologic screening | -24
no evidence of extracardiac disease | -24
cardiac magnetic resonance imaging | -24
tumourous myocardial isointense mass | -24
diffuse infiltration of the myocardium | -24
extension into the pericardium | -24
infiltration of tricuspid valve insertion | -24
referred to cardiac surgery centres | -168
deemed inoperable | -168
active surveillance | -168
best supportive therapy | -168
presentation with fatigue and dizziness | -72
atrioventricular block II type Mobitz II | -72
massive progression of the tumour mass | -72
subtotal obstruction of the tricuspid valve | -72
infiltration of the cardiac base | -72
infiltration of the atrial septum | -72
transpericardial infiltration of the diaphragm | -72
bilateral axillary lymph nodes | -72
enlargement of lymph nodes | -72
epicardial right ventricle single lead pacemaker | -72
lymph node excision | -72
histological proof of diffuse large B-cell non-Hodgkin-lymphoma | -72
pre-phase treatment with rituximab and prednisolone | -72
reduced-dose chemotherapy | -72
R-mini-CHOP | -72
continuation of chemotherapy | 0
five cycles of R-CHOP | 24
complete remission | 168
no remaining cardiac mass | 168
no extracardiac disease | 168
no AV conduction disorder | 168
18-fluorine-flurodeoxyglucose positron tomography/computed tomography | 168
pacemaker showed no stimulation | 168
no arrhythmia burden | 168