40 years old | 0
male | 0
tricuspid atresia | -25200
post-lateral tunnel Fontan | -25200
HIV | -4032
gout | 0
obstructive sleep apnea | 0
fever | -72
shortness of breath | -72
diarrhea | -72
nasopharyngeal swab test result positive for SARS-CoV-2 | -72
worsening shortness of breath | 0
presentation to the emergency department | 0
heart rate of 118 beats/min | 0
blood pressure of 159/100 mm Hg | 0
respiratory rate of 50 breaths/min | 0
oxygen saturation of 40% on room air | 0
oxygen saturation of 86% with high-flow nasal cannula | 0
left-sided pneumothorax | 0
chest x-ray film | 0
ectopic atrial rhythm/tachycardia | 0
right bundle branch block | 0
QRS duration of 113 ms | 0
QTc interval of 480 ms | 0
ejection fraction of 25% to 35% | -10080
severe aortic regurgitation | -10080
mild mitral valve regurgitation | -10080
sinus rhythm with evidence of wandering atrial pacemaker | -10080
isolated premature atrial contractions | -10080
losartan | -10080
allopurinol | -10080
ergocalciferol | -10080
elvitegravir-cobicistat-emtricitabine-tenofovir-alafenamide | -10080
normal CD4 count | -10080
pneumonia | 0
pulmonary edema | 0
atelectasis | 0
pulmonary arteriovenous malformations | 0
anemia | 0
depressed ventricular function | 0
atrioventricular valve regurgitation | 0
tamponade | 0
sepsis | 0
venovenous collaterals | 0
Fontan baffle leak | 0
increased pulmonary vascular resistance | 0
restrictive atrial communication | 0
pulmonary venous hypertension | 0
pulmonary artery obstruction | 0
large left pneumothorax | 0
collapse of the left upper and middle lung lobes | 0
abnormal laboratory test values | 0
white blood cell count of 8,000/μl | 0
hemoglobin of 15.8 g/dl | 0
hematocrit of 48% | 0
platelets of 182,000/μl | 0
sodium of 133 mmol/l | 0
chloride of 92 mmol/l | 0
aspartate transaminase of 92 U/l | 0
alanine aminotransferase of 43 U/l | 0
ferritin of 1,318 ng/ml | 0
lactate dehydrogenase of 770 U/l | 0
D-dimer of 1.37 μg/ml | 0
fibrinogen of 592 mg/dl | 0
N-terminal pro-brain natriuretic peptide of 248 pg/ml | 0
CD4 count of 142 /μl | 0
pigtail chest tube placement | 0
high-flow nasal cannula at 30 L and 100% fraction of inspired oxygen | 0
nitric oxide at 40 parts per million | 0
solumedrol 32 mg daily for 10 days | 0
remdesivir 100 mg daily for 5 days | 0
convalescent plasma | 0
transfer from the intensive care unit to the floor | 192
chest tube placed to water seal | 264
decreased hemoglobin level | 264
replacement of chest tube | 264
administration of 2 U of packed red cells | 264
nasal cannula oxygen support weaned to 1 liter | 264
discharge | 480
fatigued | 528
oxygen saturation on room air returned to baseline at rest | 528
desaturation with activity | 528