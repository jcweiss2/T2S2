3562 grams | 0
    male | 0
    admitted to the hospital | 0
    severe respiratory distress | 0
    meconium aspiration syndrome | 0
    perinatal depression | 0
    suspected neonatal sepsis | 0
    intubation | 0
    ventilator support | 0
    surfactant meconium lavage | 0
    surfactant replacement therapy | 0
    antibiotics for neonatal sepsis prophylaxis | 0
    ampicillin | 0
    gentamicin | 0
    umbilical venous catheter placement | 0
    umbilical arterial catheter placement | 0
    negative blood workup for sepsis | 0
    improving respiratory status | 0
    hypoxia resolving | 0
    respiratory acidosis resolving | 0
    weaned to minimal ventilator settings | 144
    preparation for extubation | 144
    liver enlargement noted on abdominal X-ray | 144
    mildly elevated liver enzymes | 144
    febrile | 144
    hemodynamically stable | 144
    presumptive diagnosis of disseminated neonatal HSV infection | 144
    acyclovir started | 144
    HSV polymerase chain reaction pending | 144
    blood culture repeated | 144
    blood cell parameters repeated | 144
    ampicillin continued | 144
    gentamicin continued | 144
    endotracheal tube removed | 168
    extubated to nasal cannula | 168
    failed extubation due to upper airway edema | 174
    failure of extubation due to worsening respiratory status | 174
    progressively increased abdominal girth | 174
    moderately high liver enzymes | 180
    paucity of bowel gas on chest X-ray | 180
    UVC tip at T10 | 180
    UVC migrated into the liver | 180
    insidious onset of abdominal distension | 180
    ascites | 180
    liver enlargement | 180
    markedly elevated liver enzymes | 180
    obstructive uropathy | 180
    progressive worsening of respiratory status | 180
    abdominal girth increased by 5 cm | 192
    liver size increased | 192
    chest and abdomen X-ray showing small lung volume | 192
    compressed by gasless abdomen | 192
    huge liver | 192
    marked abdominal distension | 192
    ascites | 192
    aspartate transaminase increased from 173 to 929 U/L | 192
    alanine transaminase increased from 82 to 380 U/L | 192
    total bilirubin increased from 2.7 to 4.1 g/dL | 192
    direct bilirubin increased from previous day | 192
    lactate dehydrogenase 1861 IU/L | 192
    abdominal ultrasound confirmed ascites | 192
    echogenic mass within liver | 192
    mild left hydroureter | 192
    hydronephrosis | 192
    obstructive uropathy | 192
    intrahepatic biliary duct dilatation | 192
    TPN extravasation via UVC suspected | 192
    UVC infusion stopped | 192
    UVC removed | 192
    peripheral IV access obtained | 192
    dextrose with electrolytes started | 192
    pediatric surgeon consulted | 192
    exploratory laparotomy performed | 192
    clot removal | 192
    ascites drainage | 192
    Penrose drain placement | 192
    paracentesis confirmed TPN extravasation | 192
    peritoneal fluid analysis showed protein 1213 mg/dL | 192
    peritoneal fluid analysis showed triglyceride 591 mg/dL | 192
    peritoneal fluid analysis showed glucose 539 mg/dL | 192
    HSV polymerase chain reaction negative | 240
    IV acyclovir discontinued | 240
    repeat blood culture negative | 240
    IV ampicillin discontinued | 264
    IV gentamicin discontinued | 264
    clinical status improved significantly | 240
    ascites drained | 192
    peritoneal blood clots removed | 192
    Penrose drain removed after 5 days | 336
    two 20 mL/kg packed red blood cell transfusions | 192
    anemia due to liver laceration | 192
    anemia due to hemorrhage | 192
    elevated liver enzymes normalized | 336
    hematuria resolved | 336
    enteric nutrition started | 288
    full enteric feedings attained | 456
    extubated to room air | 456
    nipple feeding started | 600
    breast feeding started | 600
    bottle feeding started | 600
    Similac Advance started | 600
    liver laceration resolved | 672
    liver mass resolved | 672
    obstructive uropathy resolved | 672
    ascites resolved | 672
    normal liver function tests | 672
    normal renal function tests | 672
    abdominal ultrasound normal | 648
    small residual liver mass | 648
    discharge home | 672