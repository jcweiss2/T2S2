26 years old | 0
male | 0
admitted to the hospital | 0
frank haematuria | -720
colicky abdominal pain | -720
increased urinary frequency | -720
dysuria | -720
treated for urinary tract infection | -720
CT abdomen demonstrated moderate bilateral hydronephrosis | -720
no calculi | -720
Common bile duct (CBD) was measured at 8 mm | -720
cystoscopy revealed a diffusely inflamed bladder | -720
marked reduction in capacity (150 cc) | -720
no obstruction at the ureteric orifices | -720
bladder biopsy showed inflammatory change | -720
no dysplasia or malignancy | -720
discharged with outpatient follow-up | -720
increasing flank pain | -96
became drowsy | -96
short of breath | -96
low blood pressure | 0
tachycardia | 0
tachypnoea | 0
Glasgow coma scale was 13/15 | 0
no localizing neurological signs | 0
severe metabolic acidosis | 0
acute renal failure | 0
abnormal liver function tests | 0
obstructive pattern | 0
regular user of street ketamine | -168
deteriorated quickly | 1
worsening respiratory function | 1
requiring intubation | 1
bilateral basal consolidation | 1
aspiration | 1
transferred to the intensive care unit | 1
vasopressors were required | 1
continuous haemofiltration (CVVH) | 1
broad-spectrum antibiotics | 1
blood cultures grew methicillin-sensitive staphylococcus aureus | 2
repeat renal ultrasound confirmed hydronephrosis | 2
bilateral nephrostomies were placed | 2
gelatinous debris was aspirated | 2
ketamine metabolites | 2
cannabanoids | 2
lignocaine | 2
dilated CBD | 2
urine output began to return | 48
bilateral nephrostograms showed free flow of contrast | 48
CVVH then intermittent dialysis | 48
renal function began to recover | 576
nephrostomies were clamped | 576
nephrostomies were removed | 576
serum creatinine was 123 μmol/l | 576
hydronephrosis had completely resolved | 576
liver function tests improved | 576
CBD dilatation resolved | 576
readmitted | 1008
right upper quadrant pain | 1008
marked derangement of liver function tests | 1008
biliary dilatation had recurred | 1008
renal tract appeared normal | 1008
serum creatinine had risen | 1008
urine analysis was positive for ketamine metabolites | 1008
treated for biliary sepsis | 1008
improvement of symptoms | 1010
underwent endoscopic retrograde cholangiopancreatography (ERCP) | 1010
no strictures or stones were seen in the CBD | 1010
stent was placed | 1010
developed pancreatitis | 1012
liver function tests had only partially improved | 1344
serum creatinine had risen | 1344
renal biopsy was performed | 1344
tubular injury and regeneration | 1344
normal vasculature and interstitium | 1344
acute tubular necrosis | 1344
sepsis and pancreatitis | 1344