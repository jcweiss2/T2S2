male | 0 | 0 | Factual
25 years old | 0 | 0 | Factual
primigravida | 0 | 0 | Factual
uncomplicated pregnancy | -280 | 0 | Factual
spontaneous onset of labor | -1 | 0 | Factual
fetal distress | -1 | 0 | Factual
ventouse-assisted delivery | 0 | 0 | Factual
birth weight 3940 grams | 0 | 0 | Factual
resuscitation with mask ventilation | 0 | 0 | Factual
intubated | 0.13 | 0.13 | Factual
transferred to NICU | 0.13 | 0.13 | Factual
synchronized intermittent positive pressure ventilation (SIPPV) | 0.13 | 13.5 | Factual
gentamicin | 0 | 120 | Factual
benzyl penicillin | 0 | 120 | Factual
neutropenia | 18 | 18 | Factual
elevated inflammatory markers | 18 | 18 | Factual
C-reactive protein (CRP) 60 mg/L | 18 | 18 | Factual
procalcitonin 68.55 µg/L | 18 | 18 | Factual
lumbar puncture | 23 | 23 | Factual
normal cell count | 23 | 23 | Factual
negative for pathogens | 23 | 23 | Factual
placental surface eSwab | 23 | 23 | Factual
Gram-negative diplococci | 23 | 23 | Factual
Neisseria meningitidis | 23 | 23 | Factual
molecular testing | 23 | 23 | Factual
N. meningitidis genogroup W | 23 | 23 | Factual
clonal complex 11 (CC11) | 23 | 23 | Factual
blood cultures negative | 0.48 | 0.48 | Factual
heel-prick blood in EDTA | 5.5 | 5.5 | Factual
N. meningitidis genogroup W DNA | 5.5 | 5.5 | Factual
benzylpenicillin dosage decreased | 13.5 | 13.5 | Factual
cefotaxime | 13.5 | 120 | Factual
maternal bloods taken | -2.5 | -2.5 | Factual
elevated leucocyte count | -2.5 | -2.5 | Factual
neutrophil count | -2.5 | -2.5 | Factual
mother remained well | 0 | 192 | Factual
baby discharged | 192 | 192 | Factual
contact tracing | 192 | 192 | Factual
chemoprophylaxis with ciprofloxacin | 192 | 192 | Factual
quadrivalent conjugate meningococcal vaccine | 192 | 192 | Factual
counseling | 192 | 192 | Factual
funisitis | -1 | 0 | Factual
chorioamnionitis | -1 | 0 | Factual
maternal and fetal inflammatory response | -1 | 0 | Factual
early-onset neonatal sepsis | 0 | 192 | Factual
invasive meningococcal disease (IMD) | 0 | 192 | Factual
N. meningitidis W CC11 | 0 | 192 | Factual