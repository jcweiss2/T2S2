63 years old | 0\
female | 0\
splenectomy | -77424\
idiopathic thrombocytopenic purpura | -77424\
menometrorhagia | -77424\
vaccinated with PPV23 | -120\
general body malaise | -48\
diarrhea | -48\
vomiting | -48\
influenza-like symptoms | -48\
confused | 0\
fever | 0\
hypotension | 0\
bradycardia | 0\
tachypnea | 0\
decreased oxygen saturation | 0\
cyanosis | 0\
severe sepsis | 0\
volume therapy | 0\
broad-spectrum antimicrobial therapy | 0\
hydrocortisone | 0\
white blood cell count | 0\
neutrophils | 0\
hemoglobin | 0\
thrombocytes | 0\
C-reactive protein | 0\
P-lactate | 0\
aB-P-O2 | 0\
aB-P-CO2 | 0\
aB-pH | 0\
Streptococcus pneumococcal urinary antigen test | 0\
discrete pulmonic stasis | 0\
disseminated intravascular coagulation | 24\
microthrombi | 24\
growth of S. pneumoniae | 48\
antimicrobial treatment changed to penicillin G | 48\
suspicion of endocarditis | 72\
modest hypokinesia of the apical part of the left ventricle | 72\
ejection fraction of 45% | 72\
endocarditis dismissed | 72\
necrosis of the fingertips and toes | 72\
renal insufficiency | 72\
hemodialysis | 72\
antibiotic therapy altered to ceftriaxone | 72\
leucocytes decreased | 96\
CRP decreased | 96\
fever dissolved | 96\
tracheal secret for culture | 96\
culture negative | 96\
transferred from the ICU to the medical department | 216\
antibiotics stopped | 216\
serological analysis of the pneumococcal isolate | 216\
serotype 12F | 216\
discharged | 528\
oral dicloxacillin | 528\
raised leucocytes | 528\
CRP | 528\
necrotic tissue on fingers and toes | 528\
wound cultures | 528\
Staphylococcus aureus | 528\
haemolytic streptococci group C/G | 528\
new TTE | 528\
amputated | 912\
readmitted with severe sepsis | 1512\
sepsis regimen | 1512\
ceftriaxone therapy | 1512\
transesophageal echocardiography | 1512\
endocarditis | 1512\
antimicrobial treatment altered to penicillin G | 1512\
treated conservatively with penicillin G | 1512\
recovered | 1596\
serological tests of the pneumococcal capsule polysaccharides | 1596\
serotype 12F | 1596\
antibodies to 12F | 1596\
antibody response to serotype 12F | 1596