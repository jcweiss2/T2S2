63 years old | 0
female | 0
admitted to the hospital | 0
fever | -48
chills | -48
malaise | -48
cigarette smoking | -6720
breast cancer resection | -6720
dog hand bite | -48
creatinine 1.22 mg/dl | 0
lactate dehydrogenase (LDH) 298 | 0
AST 115 | 0
ALT 54 U/l | 0
hyponatremia 130 mmol/l | 0
hyposmolality 265 mOsm/kg | 0
PaO2/FiO2 ratio (P/F) 246 mmHg | 0
bilateral basal hyperdensities of the lungs | 0
thrombocytopenia | 24
acute kidney injury (AKI) | 24
livedo reticularis | 24
arterial hypotension | 24
acute hypoxemic respiratory failure | 24
high serum procalcitonin (79.7 ng/ml) | 24
Gram staining of the blood culture showed thin and slender Gram-negative rods | 24
meropenem | 24
intubated | 24
septic shock (SOFA 21) | 24
severe lactic acidosis (pH 6.7, lactate 17 mmol/l) | 24
high-dose inotropic support (norepinephrine 0.5–1 μg/kg/min) | 24
continuous mandatory mechanical ventilation (P/F 90) | 24
hydrocortisone 200 mg/die | 24
renal replacement therapy using continuous venovenous hemodialysis (CVVHD) | 72
rhabdomyolysis | 96
liver injury | 96
severe thrombocytopenia | 96
coagulopathy | 96
fresh frozen plasma and platelet transfusion | 96
livedo reticularis worsened to a frank purpura | 96
ischemia of the limbs | 96
ampicillin-sulbactam and ceftriaxone | 168
surgical amputation of her finger | 336
end-stage renal disease | 5760
intermittent hemodialysis | 5760