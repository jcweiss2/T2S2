28 years old | 0
female | 0
admitted to the hospital | 0
twin pregnancy | 0
Sheehan syndrome | 0
gravida 2 | 0
live 0 | 0
pyrexia | -720
pyonephritis | -720
severe hyperglycemia | -720
metabolic acidosis | -720
septicemic shock | -720
bilateral pleural effusion | -720
respiratory distress | -720
loss of fetus | -720
drainage of pus | -720
broad-spectrum antibiotics | -720
hemodialysis | -720
hypothyroidism | -624
equivocal serum cortisol levels | -624
pituitary apoplexy | -624
hydrocortisone | -624
thyroxine | -624
intrauterine insemination | -624
conceived | -624
diamniotic monochorionic twins | -624
gestational diabetes mellitus | -624
elective lower segment cesarean section | 0
multiple metabolic derangements | 0
intrauterine growth retardation | 0
subarachnoid block | 0
invasive blood pressure monitoring | 0
perioperative intravenous hydrocortisone supplementation | 0
nil per oral | -8
thyroxine | -2
ranitidine | -2
metoclopramide | -2
fasting blood sugar | -2
insulin withheld | -2
hydrocortisone | 0
electrocardiogram | 0
pulse oximetry | 0
noninvasive blood pressure monitoring | 0
wide bore i/v cannulae | 0
arterial cannula | 0
supplemental oxygen | 0
subarachnoid block administered | 0
bupivacaine | 0
fentanyl | 0
surgery commenced | 0
hypotension | 6
phenylephrine | 6
live male babies | 60
APGAR scores | 60
oxytocin infusion | 60
intraoperative blood loss | 60
surgery duration | 60
intraoperative arterial blood gas analysis | 60
postoperative pain relief | 120
paracetamol | 120
high dependency unit | 120
postoperative period | 168
follow-up | 168
discharged | 168