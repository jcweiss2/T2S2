52 years old | 0
male | 0
admitted to the hospital emergency room | 0
general weakness starting | -240
right upper quadrant pain | -96
PC-type MCD diagnosed | -43800
multiple lymph node enlargements in neck, axillary, mediastinal, abdominal, and pelvic space | -43800
right axillary lymph node biopsy under local anesthesia | -43800
eight cycles of chemotherapy | -43800
complete remission | -43800
loss to follow-up | -43800
no history of taking specific drugs | -43800
smoking history of 20 pack-years | -43800
acute calculous cholecystitis | 0
lymphadenopathy with multiple enlarged nodes in abdomen and pelvis | 0
splenomegaly | 0
bilateral pleural effusion | 0
small amounts of ascites in cul-de-sac | 0
anemia | 0
thrombocytopenia | 0
lymphopenia | 0
azotemia | 0
stress-induced cardiomyopathy (EF=43%) | 0
percutaneous transhepatic gallbladder drainage | 0
multiple lymph node enlargements | 0
suspicion of recurrence of CD | 0
evaluation | 0
polyclonal hypergammaglobulinemia | 0
plasmacytosis | 0
reductions in platelet count | 0
reductions in hemoglobin | 0
reductions in lymphocyte | 0
reductions in total cholesterol | 0
reductions in albumin | 0
increases in INR | 0
increases in blood urea nitrogen | 0
increases in creatinine | 0
increases in CRP | 0
increases in ESR | 0
increases in VEGF | 0
serological test for HIV negative | 0
started on chemotherapy | 0
pulmonary edema worsened | 168
stress-induced cardiomyopathy exacerbation (EF=25%) | 168
dyspnea | 168
oliguria | 168
aggressive treatment including ICU admission | 168
clinical signs gradually improved | 168
normalization of left ventricular systolic function (EF=68%) | 552
improvements in pulmonary edema | 552
improvements in azotemia | 552
transfusions of leukocyte-poor and irradiated packed RBC | 552
transfusions of platelets | 552
transfusions of FFP | 552
no significant improvement in blood lab values | 552
Hgb 3.8-11.6 g/dl | 552
platelet count 31,000-132,000/µl | 552
INR 1.32-2.02 | 552
elective laparoscopic cholecystectomy planned | 720
preanesthetic evaluation performed | 720
blood transfusion of 2 units RBC | 720
blood transfusion of 8 units platelets | 720
blood transfusion of 4 units FFP | 720
Hgb 9.0 g/dl | 720
platelet 78,000/µl | 720
INR 1.41 | 720
mild dyspnea | 720
no cough | 720
no sputum | 720
abdominal distension | 720
chest X-ray showing ill-defined consolidation in both lungs | 720
no rales | 720
no wheezing | 720
pulmonary function test not performed | 720
ECG normal | 720
thoracic CT scan no mediastinal mass | 720
transferred to operating room | 720
ECG monitoring | 720
pulse oximetry monitoring | 720
bispectral index monitoring | 720
modified Allen's test performed | 720
22 G catheter inserted in left radial artery | 720
FloTrac/Vigileo monitor connected | 720
room air ABGA: pH 7.53 | 720
room air ABGA: PaCO2 27 mmHg | 720
room air ABGA: PaO2 65 mmHg | 720
room air ABGA: HCO3- 22.6 mEq/L | 720
room air ABGA: BE -0.1 mEq/L | 720
room air ABGA: SaO2 95% | 720
room air ABGA: Hgb 8.8 g/dl | 720
room air ABGA: Hct 26% | 720
electrolytes normal | 720
general anesthesia induced | 720
intravenous thiopental sodium 100 mg | 720
intravenous lidocaine 40 mg | 720
intravenous etomidate 10 mg | 720
intravenous cisatracurium 14 mg | 720
intravenous remifentanil 0.15 µg/kg/min | 720
tracheal tube inserted orotracheally | 720
general anesthesia maintained with sevoflurane 1.5-3 vol% | 720
O2 1.5 L/min | 720
air 1.5 L/min | 720
remifentanil 0.05 µg/kg/min | 720
PreSep central venous oximetry catheter inserted via right internal jugular vein | 720
foley catheter not inserted | 720
Vigileo monitor parameters monitored | 720
Calot's triangle severe inflammation and adhesion | 720
dissection impossible | 720
surgery switched to open cholecystectomy | 720
perioperative drainage of ascites 2 L | 720
additional cisatracurium 2 mg | 720
additional ephedrine 5 mg | 720
BP 105-150/50-85 mmHg | 720
HR 82B110 beats/min | 720
oxygen saturation 100% | 720
Vigileo parameters normal | 720
bispectral index 32-39 | 720
ABGA during surgery: pH 7.39 | 720
ABGA during surgery: PaCO2 38 mmHg | 720
ABGA during surgery: PaO2 141 mmHg | 720
ABGA during surgery: HCO3- 23 mEq/L | 720
ABGA during surgery: BE -2 mEq/L | 720
ABGA during surgery: SaO2 99% | 720
ABGA during surgery: Hgb 7.8 g/dl | 720
ABGA during surgery: Hct 23% | 720
ABGA during surgery: Na 138 mmol/L | 720
ABGA during surgery: K 3.8 mmol/L | 720
ABGA during surgery: Ca2+ 0.97 mmol/L | 720
surgery uneventful | 720
operation duration 1.5 hours | 720
anesthesia duration 2.5 hours | 720
no significant blood loss | 720
infused crystalloid fluid 1,100 ml | 720
anesthesia terminated | 720
patient awakened smoothly | 720
tracheal tube removed | 720
transferred to ICU | 720
postoperative vital signs satisfactory | 720
postoperative laboratory findings satisfactory | 720
moved to general ward next day | 768
continuous chemotherapy for CD | 768
cough developed | 1440
sputum developed | 1440
fungal pneumonia suspected | 1440
treatment started | 1440
condition rapidly deteriorated | 1440
aggressive treatment including ventilator care in ICU | 1440
expired | 1512
