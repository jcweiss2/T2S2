49 years old | 0
    male | 0
    admitted to the hospital | 0
    spider bite on right shoulder | -120
    doxycycline prescription | -72
    worsening rash | -48
    fever | -48
    body aches | -48
    discoloration of urine | -48
    sepsis criteria met | -48
    refusal of hospital admission | -48
    pain around bite | -24
    chest pain | -24
    fevers | -24
    body aches | -24
    shortness of breath | -24
    nausea | -24
    vomiting | -24
    black colored urine | -24
    hemolysis | 0
    acute renal failure | 0
    intravenous vancomycin | 0
    piperacillin/tazobactam | 0
    admission to intensive care unit | 0
    hemodialysis recommendation | 0
    antibiotics de-escalation | 0
    supportive care for spider bite | 0
    packed red blood cell transfusion | 0
    hemoglobin/hematocrit monitoring | 0
    acute hemolytic anemia | 0
    no thrombotic microangiopathy | 0
    complement-mediated hemolysis | 0
    worsening acute kidney injury | 48
    nausea | 48
    vomiting | 48
    oliguria | 48
    hemodialysis line placement | 48
    intermittent hemodialysis | 48
    additional packed red blood cell transfusion | 48
    plasmapheresis initiation | 72
    albumin replacement | 72
    packed red blood cell transfusion post-plasmapheresis | 72
    antibiotics broadening | 72
    ultrasound of spider bite site | 72
    second plasmapheresis | 120
    clinical improvement | 120
    folic acid initiation | 120
    three hemodialysis sessions | 120
    discharge | 168
    close follow-up | 168
    outpatient labs | 168
    creatinine improvement | 168
    white blood cell count improvement | 168
    hemoglobin improvement | 168
    platelet count improvement | 168
    
