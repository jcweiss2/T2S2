30 years old | 0
female | 0
history of polysubstance abuse | 0
anxiety | 0
depression | 0
unresponsive | 0
found in a bathtub | -1
injected intravenous heroin | -1
NARCAN administered | -1
no improvement of respiratory status | -1
no improvement of level of consciousness | -1
arrived at ED | 0
did not respond to verbal or painful stimuli | 0
intermittently moaning | 0
NARCAN administered intravenously | 0
no significant improvement in mental status | 0
intubated | 0
etomidate administered | 0
succinylcholine administered | 0
axillary temperature 25.8°C | 0
pulse rate 55 | 0
respiratory rate 16 | 0
blood pressure 94/40 | 0
wet clothes removed | 0
warm blankets applied | 0
temperature-sensing Foley inserted | 0
clear yellow urine returned | 0
topical warming with Bair Hugger system | 0
warm saline bags applied | 0
warmed IV normal saline administered | 0
hyperkalemia | 0
creatinine 1.16 mg/dL | 0
hyperglycemia | 0
hypocalcemia | 0
leukocytosis | 0
atrial fibrillation | 0
Osborne waves | 0
central venous access obtained | 1
transferred to intensive care unit | 1
warm IV fluids administered | 1
bladder irrigation | 1
insulin administered | 1
calcium gluconate administered | 1
normotensive | 2
normothermic | 2
repeat EKG obtained | 2
normal rate | 2
normal rhythm | 2
normal QRS complex | 2
Osborne waves resolved | 2
extubated | 24
following commands | 24
answering questions appropriately | 24
discharged home | 72
friends placed her in the bathtub | -2
friends filled the tub with ice | -2
ice cubes inserted rectally | -2