47 years old | 0
female | 0
admitted to the hospital | 0
fever | -96
left loin pain | -96
autosomal dominant polycystic kidney disease | -672
polycystic liver disease | -672
tobacco use denied | 0
alcohol use denied | 0
blood pressure 127/91 mmHg | 0
heart rate 133 beats/min | 0
respiratory rate 20/min | 0
body temperature 38.5 °C | 0
hard mass at the level of the belly button on the right abdomen | 0
no tenderness in the abdomen | 0
percussion pain in the left kidney area | 0
leukocytosis | 0
platelet count 97 × 10^9/L | 0
C-reactive protein level 214.5 mg/L | 0
serum creatinine level 97.6 μmol/L | 0
plasma fibrinogen level 6.63 g/L | 0
numerous white blood cells in the urine | 0
multiple air pockets in the left collecting system | 0
multiple hypodense cysts in bilateral kidneys | 0
multiple renal stones located in left pelvis | 0
left hydronephrosis | 0
insertion of a double “J” stent | 48
oral antibiotic treatment (nitrofurantoin 100 mg q8 h) | 0
condition rapidly deteriorated | 48
intraoperative findings revealed pus in the left collecting system | 48
culture of pus yielded ESBL positive Escherichia coli | 48
intravenous antibiotics changed to imipenem-cilastatin | 48
postoperative CT showed air spaces in the left collecting system had disappeared | 72
left hydronephrosis significantly improved | 72
discharged on day 18 | 432
readmitted 2 mo postoperatively | 1440
removal of stones from the left renal pelvis | 1470
oral antibiotic treatment (nitrofurantoin 50 mg q8 h) | 1440
flexible ureteroscopy lithotripsy | 1470
shivering 2 h postoperatively | 1472
blood pressure 60/40 mmHg | 1472
heart rate 133/min | 1472
temperature 41°C | 1472
white blood cell count significantly decreased | 1472
severe hematuria | 1472
transferred to the intensive care unit | 1472
intravenous antibiotics (meropenem 1.0 g q8 h) | 1472
right internal jugular vein punctured | 1472
norepinephrine prescribed | 1472
right radial artery punctured | 1472
600 mL of fresh plasma transfused | 1472
blood cultures performed | 1472
general condition improved | 1476
transferred back to the general ward | 1476
continued meropenem treatment | 1476
postoperative CT showed stones in the left renal pelvis had been cleared | 1500
discharged on the 23rd day | 1656
follow-up for 44 mo | 21120
serum creatinine remained below 100 μmol/L | 21120
CT showed no stones in the left renal pelvis | 21120
stones in the lower calyx significantly smaller in size and fewer in number | 21120