75 years old | 0
female | 0
habit of taking vinegar daily for 50 years | -438000
hypertension | -438000
amlodipine 10 mg daily | -438000
transported to emergency room | 0
vomiting | 0
loss of consciousness | 0
unconscious | 0
hypotensive | 0
respiratory failure | 0
blood pressure 86/58 mmHg | 0
sinus tachycardia | 0
oxygen saturation 90% | 0
no subcutaneous emphysema | 0
no signs of peritoneal irritation | 0
white blood count 3500 | 0
C-reactive protein 8.7 mg/dL | 0
renal dysfunction | 0
electrolytes within normal ranges | 0
liver function within normal ranges | 0
urinalysis within normal ranges | 0
computed tomography showed poor contrast in middle intrathoracic esophagus | 0
mediastinal emphysema | 0
right pneumothorax | 0
pleural effusion | 0
diagnosed with septic shock due to esophageal rupture | 0
emergency surgery | 0
opened chest through posterolateral incision of sixth intercostal space | 0
left-sided supine position | 0
right chest cavity highly contaminated with fluid containing food residue | 0
25 mm perforation in middle intrathoracic esophagus | 0
esophageal mucosa turned black | 0
suture closure not possible | 0
resected thoracic esophagus by 10 cm | 0
needed esophageal fistula | 0
needed enteric fistula | 0
shock vitals prolonged intraoperatively | 0
immediate systemic management in ICU | 0
esophagectomy | 0
intrathoracic lavage drainage | 0
excised specimen showed blackened esophageal mucosa | 0
no obvious malignant findings | 0
histopathological examination revealed ulcerated and necrotic esophageal mucosa | 0
perforation in one place | 0
lymphocytic infiltration in mucosal surface layer | 0
no findings beyond muscle layer | 0
cause of perforation undetermined | 0
intensive care started immediately after surgery | 24
vitals stable 15 hours postoperatively | 39
performed esophageal fistula | 39
performed enteric fistula | 39
esophageal fistula mucosa blackened | 39
esophageal fistula mucosa normalized on seventh postoperative day | 168
general condition improved sufficiently | 1440
underwent esophageal reconstruction by third operation 60 days after first operation | 1440
posterior sternal pathway cervical esophagogastric anastomosis | 1440
cholecystectomy | 1440
started oral intake on 12th day after third surgery | 360
discharged on 27th day after third surgery | 648
