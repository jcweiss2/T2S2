26 years old|0
    male|0
    admitted in the emergency department|0
    weakness of all four limbs|-24
    pharmacist at a private nursing home|0
    addicted to multiple medicines including tramadol, diclofenac, pheniramine, and dexamethasone|0
    addicted to heparin|0
    bronchial asthma|0
    on and off steroids|0
    conscious|0
    oriented|0
    hemodynamically stable|0
    heart rate of 112 beats/min|0
    non-invasive blood pressure of 130/80 mmHg|0
    respiratory rate of 24/min|0
    temperature of 99°F|0
    no pallor|0
    no signs of clubbing|0
    no lymphadenopathy|0
    oral thrush present|0
    chest examination grossly normal|0
    cardiovascular system examination grossly normal|0
    per abdomen examination grossly normal|0
    power grade 3/5 in upper limbs|0
    power grade 1/5 in lower limbs|0
    generalized areflexia|0
    planters bilateral flexors|0
    sensory examination normal|0
    arterial blood gas (ABG) at admission showed normal pH (7.437)|0
    hyperkalemia (K+ = 6.01)|0
    admitted to intensive care unit|0
    tachypnoeic|-1
    respiratory rate of 36-40/min|-1
    non-invasive ventilation|-1
    heart rate 130 beats/min|-1
    pulses feeble|-1
    blood pressure 100/56 mmHg|-1
    invasive lines|-1
    central venous cannulation|-1
    arterial line|-1
    central venous pressure 6 cm H2O|-1
    mean arterial pressure (MAP) 55 mmHg|-1
    resuscitated with 1 litre normal saline|-1
    blood pressure improved|0
    MAP 64 mmHg|0
    given 500 mL normal saline|0
    started on normal saline 100 mL/h infusion|0
    MAP of >65 mmHg targeted|0
    urine output >0.5 mL/kg|0
    chest X-ray showed patch of consolidation on the right middle and lower zones|0
    echocardiography showed global hypokinesia|0
    severe left ventricular dysfunction|0
    ejection fraction of 30%|0
    repeat ABG after 6 h showed metabolic acidosis|6
    lactic acidosis|6
    hyperkalemia (K+ = 7.0)|6
    S. K+ 6.7 mEq/L|6
    anti-hyperkalemia treatment started|6
    calcium gluconate|6
    dextrose-insulin|6
    salbutamol nebulization|6
    slow low-efficiency dialysis (SLED) of 8 h|6
    pulseless ventricular tachycardia|6.33
    defibrillated|6.33
    CPR done|6.33
    anti-hyperkalemia regimen repeated|6.33
    serum K+ 9.1 mEq/L|6.33
    revived after 40 min CPR|6.67
    intubated|6.67
    invasive ventilatory support|6.67
    started on inotropes|6.67
    started on vasopressors|6.67
    subsequent ABG showed persistent hyperkalemia (K+ = 7.1)|8
    pH improvement|8
    extended SLED|8
    SLED total duration 20 h|20
    post dialysis serum K+ 7.6 mEq/L|20
    developed blisters all over the body|20
    coagulopathy|20
    thrombocytopenia (platelets 33,000/mm3)|20
    PT/INR increased from 1.21 to 6.8|20
    sepsis suspected|20
    started on ceftriaxone|0
    shifted to meropenem|20
    shifted to teicoplanin|20
    shifted to ampicillin|20
    deterioration in blood gas showing acidosis|24
    rise in potassium levels|24
    SLED again|24
    dialyzed for more than 32 h|32
    hyperkalemia refractory to antihyperkalemic agents|40
    high anion gap acidosis|40
    fludrocortisone 100 μg/day|48
    activated clotting time monitored|48
    protamine sulphate given|48
    upper gastrointestinal bleed|72
    asystole|72
    CPR done|72
    declared dead|72
    blood cultures showed methicilin-resistant staphylococci|72
    