28 years old | 0
female | 0
8 weeks pregnant | 0
acute severe asthma | -10
short non-infective prodrome | -10
hypoxic cardiac arrest | -10
ventricular fibrillation | -10
resuscitation to sinus tachycardia | -10
endotracheal intubation | -10
therapeutically cooled to 33°C | 0
salbutamol | 0
ipratropium | 0
aminophylline | 0
hydrocortisone | 0
magnesium | 0
ketamine | 0
inhalation anesthesia with 1 MAC isoflurane | 0
severe hypercapnic acidosis | 0
neuromuscular blockade | 0
ventilation improving | 24
intravenous sedatives stopped | 48
NMB stopped | 48
generalised status myoclonus | 48
isoflurane stopped | 96
comatose | 96
absent motor response to painful stimulus | 96
preserved pupillary reflexes | 96
preserved corneal reflexes | 96
preserved cough reflexes | 96
preserved gag reflexes | 96
spontaneously breathing | 96
severe GSM | 96
refractory to three antiepileptic medications | 96
generalised periodic discharges on EEG | 96
no discernable background rhythm on EEG | 96
reversible causes of coma eliminated | 96
no agreement about neurological outcome | 192
social issues | 192
interethnic marriage | 192
pregnancy | 192
intensive social work support | 192
plasma neuron-specific enolase | 240
NSE 51 mcg/L | 240
somatosensory-evoked potential | 240
SSEP unhelpful due to myoclonus motion artefacts | 240
brain MRI | 240
bilateral basal ganglia infarction | 240
frontoparietal cortex infarction | 240
severe hypoxic encephalopathy | 240
medical consensus regarding poor prognosis | 240
extubated | 264
died | 288