67 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
hypertension | 0 | 0 | Factual
degenerative joint disease | 0 | 0 | Factual
bilateral knee replacement | -17472 | -17472 | Factual
substance abuse | 0 | 0 | Factual
trauma to face and chest wall | -24 | -24 | Factual
lightheadedness | 0 | 0 | Factual
fatigue | 0 | 0 | Factual
leukocytosis | 0 | 0 | Factual
hemoglobin of 10.2 g | 0 | 0 | Factual
venous lactic acid of 2.4 mol/l | 0 | 0 | Factual
intramuscular and subpectoral hematoma | 0 | 0 | Factual
extrapleural extension into the chest | 0 | 0 | Factual
acute right second through fifth anterior rib fractures | 0 | 0 | Factual
bilateral lower lobe bronchopneumonia | 0 | 0 | Factual
blood cultures obtained | 0 | 0 | Factual
empiric antibiotics with intravenous piperacillin–tazobactam | 0 | 48 | Factual
afebrile | 0 | 0 | Factual
hypotensive | 0 | 0 | Factual
admitted to intensive care unit | 0 | 0 | Factual
suspected septic shock | 0 | 0 | Factual
initiation of vasopressors | 0 | 0 | Factual
antibiotics broadened to intravenous vancomycin, cefepime and metronidazole | 48 | 96 | Factual
repeat blood, urine and sputum cultures obtained | 48 | 48 | Factual
blood and urine cultures resulted as negative | 96 | 96 | Factual
sputum cultures grew methicillin-resistant Staphylococcus aureus | 96 | 96 | Factual
antibiotics narrowed to intravenous vancomycin | 96 | 120 | Factual
left knee pain | 120 | 120 | Factual
notable swelling on physical exam | 120 | 120 | Factual
concern for infection of prosthetic knee joint | 120 | 120 | Factual
sterile left knee aspiration | 120 | 120 | Factual
synovial fluid was cloudy, amber colored | 120 | 120 | Factual
white blood cells of 9.28 × 103/mcL | 120 | 120 | Factual
calcium pyrophosphate crystals | 120 | 120 | Factual
complete washout and debridement of the joint with retention of the prosthesis | 144 | 144 | Factual
infected knee with purulence | 144 | 144 | Factual
cultures from the infected area obtained | 144 | 144 | Factual
antibiotic regimen transitioned to intravenous cefazolin | 168 | 168 | Factual
cultures resulted with C. bifermentans | 240 | 240 | Factual
antibiotic regimen transitioned to intravenous ampicillin–sulbactam | 240 | 336 | Factual
contrast computerized tomography scan of the abdomen | 240 | 240 | Factual
human immunodeficiency virus screening | 240 | 240 | Factual
discharged to a rehabilitation facility | 384 | 384 | Factual
referral to gastroenterology for outpatient colonoscopy | 384 | 384 | Factual
recovered full range of motion of left knee | 744 | 744 | Factual
no signs of lingering joint or systemic infection | 744 | 744 | Factual
taking Augmentin | 744 | 744 | Factual
medication adherence | 744 | 744 | Factual
had not yet opted to undergo colonoscopy | 744 | 744 | Factual