85 years old | 0
male | 0
admitted to the hospital | 0
fall at home | -72
lethargy | -72
productive cough | -72
decreased oral intake | -72
transfusion-dependent chronic myelomonocytic leukaemia type 1 | -720
type II diabetes mellitus | -720
atrial fibrillation | -720
permanent pacemaker | -720
chronic kidney disease stage III | -720
hypertension | -720
permanent suprapubic catheter | -720
neurogenic bladder | -720
benign prostatic hypertrophy | -720
restless leg syndrome | -720
duodenal ulcers | -720
hypercholesterolaemia | -720
renal calculi | -720
pyelonephritis | -720
infective endocarditis of the aortic valve | -720
non-ST elevation myocardial infarction | -720
polymyalgic rheumatoid arthritis | -720
chronic obstructive pulmonary disease | -720
irbesartan | -720
digoxin | -720
pantoprazole | -720
bisoprolol | -720
apixaban | -720
sulfasalazine | -720
pramipexole | -720
domperidone | -720
atorvastatin | -720
cholecalciferol | -720
mixed insulin | -720
paracetamol | -720
dicloxacillin | -720
low-grade fever | 0
blood pressure 131/47 mm Hg | 0
heart rate 70 bpm | 0
respiratory rate 21 | 0
oxygen saturation 93% | 0
crackles at the lung bases bilaterally | 0
massive splenomegaly | 0
acute kidney injury | 0
creatinine 325 μmol/L | 0
urea 28 mmol/L | 0
estimated glomerular filtration rate 14 mL/min/1.73 m2 | 0
serum glucose 14.2 mmol/L | 0
haemoglobin 80 g/L | 0
platelets 103×109/L | 0
white cell count 40.3×109/L | 0
neutrophils 22.91×109/L | 0
monocytes 13.43×109/L | 0
metabolic acidosis | 0
pH 7.31 | 0
bicarbonate 14 mmol/L | 0
lactate 1.3 mmol/L | 0
anion gap 21 mmol/L | 0
patchy perihilar opacification | 0
increased interstitial markings | 0
ceftriaxone | 0
doxycycline | 0
transfusion of packed red cells | 12
tachypnoea | 12
desaturation to 80% | 12
fluid overload | 12
respiratory crackles to mid-zones bilaterally | 12
poor urine output | 12
arterial blood gas | 24
pH 7.26 | 24
bicarbonate 10 mmol/L | 24
lactate 1.1 mmol/L | 24
anion gap 19 mmol/L | 24
inflammatory markers significantly raised | 24
C-reactive protein 165 mg/L | 24
WCC 80.4×109/L | 24
neutrophils 53.22×109/L | 24
lymphocytes 6.13×109/L | 24
monocytes 17.61×109/L | 24
eosinophils 1.15×109/L | 24
basophils 0.38×109/L | 24
piperacillin–tazobactam | 24
furosemide | 24
high-flow nasal prong oxygen | 24
diuresis | 48
acidosis persisted | 48
anion gap 21.3 mmol/L | 48
renal ultrasound | 48
multiple small calculi in the right kidney | 48
no evidence of obstruction or hydronephrosis | 48
urine highly positive for leukocytes | 48
Candida sp | 48
negative for eosinophils, casts, monoclonal immunoglobulin and Bence-Jones proteins | 48
pyroglutamic acidosis considered | 48
dicloxacillin and paracetamol withheld | 48
cephalexin recommended | 48
acceleration phase of leukaemia or transformation to CMML-2 | 48
spontaneous tumour lysis syndrome | 48
met two of the laboratory criteria for TLS | 48
increase in creatinine greater than or equal to 1.5 times the upper limit of normal | 48
fluconazole | 72
acidosis resolved | 168
bicarbonate improved to 26 mmol/L | 168
anion gap 14.8 | 168
renal function stabilised | 168
GFR 16 mL/min/1.73 m2 | 168
creatinine 292 μmol/L | 168
blood count differential stabilised | 168
WCC 20.1×109/L | 168
neutrophils 11.28×109/L | 168
monocytes 5.84×109/L | 168
basophils 0.20×109/L | 168
pyroglutamic acid levels 62 μmol/L | 168
discharged to a residential aged care facility | 240
symptomatic management and palliative care | 240