10 weeks old | 0
male | 0
admitted to the hospital | 0
severe abdominal distention | 0
lethargy | 0
fever | -72
poor feeding | -72
vomiting | -72
cessation of bowel movements | -24
progressive abdominal distention | -24
irritability | -24
lethargy | -24
born at term by vaginal delivery | -840
weight of 1.860 grams | -840
small for gestational age | -840
no delay in passing meconium at birth | -840
no history of constipation | -840
being breast fed | -840
vaccination schedule up to date | -840
no family history of Hirschsprung's disease | -840
no congenital disorders | -840
physical examination | 0
afebrile | 0
fair heart rate | 0
tachypneic | 0
hypotensive | 0
oxygen saturation on room air of 97% | 0
unwell | 0
lethargic | 0
dehydrated | 0
distended abdomen | 0
tense abdomen | 0
tender to palpation | 0
reduced bowel sounds | 0
laboratory investigations | 0
high leukocyte count | 0
neutrophilia | 0
thrombocytosis | 0
elevated C-reactive protein | 0
electrolyte disturbance | 0
hypo natremia | 0
hyperglycemia | 0
elevated liver function tests | 0
compensated metabolic acidosis | 0
plain abdominal X-ray | 0
multiple air fluid levels | 0
no pneumoperitoneum | 0
treated for clinical sepsis | 0
fluid resuscitation | 0
initiation of broad spectrum parenteral antibiotics | 0
diagnosis of complicated intestinal obstruction | 0
urgent laparotomy | 0
ileum massively dilated | 0
identification of a distal segment perforation | 0
primary repair of the ileal perforation | 0
totally collapsed microcolon | 0
transition zone identified at the ileocecal valve | 0
full thickness biopsies | 0
appendectomy | 0
protective ileostomy | 0
histological evidence of enterocolitis | 0
cardio-pulmonary arrest | 8
resuscitation | 8
cardio-pulmonary arrest | 20
resuscitation | 20
death | 20
autopsy not performed | 20
final diagnosis | 20
ileal perforation | 0
enterocolitis | 0
sepsis | 0
septic shock | 0
total colonic aganglionosis | 0
Hirschsprung's disease | 0