22 years old | 0
male | 0
temporal lobe epilepsy | -0
mental retardation | -0
sodium valproate | -0
Levetiracetam | -0
admitted to the emergency room | 0
generalized tonic clonic seizure | 0
sedated | 0
intubated | 0
admitted to the Intensive Care Unit (ICU) | 0
status epilepticus | 0
fever | 48
increased tracheobronchial secretions | 48
leukocyte count of 18.3 x 10^9/mL | 48
culture of tracheobronchial secretions showed growth of Pseudomonas aeruginosa | 48
chest X-ray showed new infiltrates in right lower lobe consolidation | 48
diagnosis of VAP | 48
extubated | 96
transferred to a ward | 120
febrile | 168
hypotensive | 168
transferred back to ICU | 168
antibiotics modified to a combination of Piperacillin-Tazobactam and Vancomycin | 168
improved clinically | 192
transferred out of ICU to ward | 192
vital signs were stable | 192
afebrile | 192
maintaining oxygen saturation on room air | 192
returned to baseline condition | 192
progressive bulbar weakness | 312
ataxia | 312
ophthalmoplegia | 312
finger to nose dysmetria | 312
dysdiadochokinesia | 312
abnormal heel to shin test | 312
generalized areflexia | 312
difficulty in standing | 312
lumbar puncture | 312
CSF analysis showed proteins 100mg/dl | 312
white cell count of 10 | 312
MRI brain and spine | 312
re-demonstration of atrophic left hippocampus | 312
abnormal T2 and Flair hyperintense signals | 312
mesial temporal sclerosis | 312
levels of anti-ganglioside antibodies were: Anti-GD1b 198, Anti-GD1a 175, Anti-GM1 154, Anti-GM2 41 and Anti-GQ1b <30 | 312
diagnosis of sero-negative MFS variant of GBS | 312
received 5 sessions of intravenous immunoglobulin (IVIG) | 315
hemodynamic status improved | 318
blood pressure reading of 113/67mmHg | 318
heart rate was 68–75 beats per minutes | 318
neurologic symptoms did not improve | 318
hemodynamic status stabilized | 318
rehabilitation team was consulted | 318
discharged | 336