38 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
13th week of pregnancy | 0 | 0 | Factual
abdominal discomfort | -24 | 0 | Factual
nausea | -24 | 0 | Factual
vomiting | -24 | 0 | Factual
no fever | -24 | 0 | Negated
no vaginal discharge | -24 | 0 | Negated
evaluated in the Obstetric Emergency Department | -24 | -24 | Factual
discharged home | -24 | -24 | Factual
persistent abdominal pain | -144 | 0 | Factual
nausea | -144 | 0 | Factual
vomiting | -144 | 0 | Factual
tachycardic | 0 | 0 | Factual
diffuse abdominal pain | 0 | 0 | Factual
guarding on the right quadrants | 0 | 0 | Factual
neutrophilia | 0 | 0 | Factual
low prothrombinemia | 0 | 0 | Factual
acute renal failure | 0 | 0 | Factual
high procalcitonin | 0 | 0 | Factual
high c-reactive protein | 0 | 0 | Factual
abdominal ultrasound | 0 | 0 | Factual
moderate fluid in all quadrants | 0 | 0 | Factual
good foetal vitality | 0 | 0 | Factual
hypotension | 0 | 0 | Factual
general abdominal guarding | 0 | 0 | Factual
hyperlacticaemia | 0 | 0 | Factual
hypokalaemia | 0 | 0 | Factual
hyperglycaemia | 0 | 0 | Factual
septic shock with an abdominal source | 0 | 0 | Factual
emergency exploratory laparotomy | 0 | 0 | Factual
generalised purulent peritonitis | 0 | 0 | Factual
perforated acute appendicitis | 0 | 0 | Factual
appendicectomy | 0 | 0 | Factual
thorough abdominal washing | 0 | 0 | Factual
laparostomy | 0 | 0 | Factual
admitted to the Intensive Care Unit | 0 | 0 | Factual
septic shock | 0 | 48 | Factual
need for vasopressor therapy | 0 | 48 | Factual
dialysis | 0 | 48 | Factual
intravenous piperacillin-tazobactam antibiotherapy | 0 | 48 | Factual
laparostomy revision | 48 | 48 | Factual
marked bowel oedema and distention | 48 | 48 | Factual
mild intraabdominal soiling | 48 | 48 | Factual
further peritoneal lavage | 48 | 48 | Factual
new laparostomy with progressive closure technique | 48 | 48 | Factual
recovered progressively | 48 | 96 | Factual
surgical revision | 96 | 96 | Factual
abdominal cavity primary closed | 96 | 96 | Factual
antibiotherapy adjusted | 144 | 144 | Factual
piperacillin-tazobactam suspended | 144 | 144 | Factual
amoxicillin with clavulanic acid started | 144 | 144 | Factual
transferred to the obstetrics ward | 288 | 288 | Factual
good foetal viability | 288 | 336 | Factual
discharged home | 336 | 336 | Factual
elective caesarean section | 1008 | 1008 | Factual
gave birth to a healthy child | 1008 | 1008 | Factual
ventral hernia | 7776 | 7776 | Factual
incisional hernia | 7776 | 7776 | Factual
child thriving without neurological or other impairments | 7776 | 7776 | Factual