42 years old | 0
    male | 0
    presented with fever | 0
    presented with cough | 0
    presented with dyspnoea | 0
    presented with headache | 0
    diagnosed with COVID-19 | 0
    RT-PCR positive for SARS-CoV-2 | 0
    physical examination | 0
    moderate systolic hypertension (155/85 mmHg) | 0
    heart rate 94 b.p.m. | 0
    respiratory rate 30 breaths/min | 0
    oxygen flow rate 15 L/min | 0
    O2 saturation 94% | 0
    use of non-rebreather mask | 0
    no signs of left ventricular failure | 0
    no leg oedema | 0
    fine scattered crackles present | 0
    electrocardiogram (ECG) normal | 0
    echocardiogram normal | 0
    chest X-ray bilateral peripheral pulmonary infiltrates | 0
    white cell count 19.5 × 10^9/L | 0
    neutrophil count 14.5 × 10^9/L | 0
    lymphocyte count 0.7 × 10^9/L | 0
    platelet count 360 × 10^9/L | 0
    haematocrit 24.6% | 0
    ferritin level 855 μg/L | 0
    high-sensitivity C-reactive protein level 112.0 mg/L | 0
    D-dimer level 4400 ng/mL | 0
    fibrinogen level 7.1 g/L | 0
    prothrombin time 17.0 s | 0
    activated partial thromboplastin time (aPTT) 43.7 s | 0
    initial treatment with ceftriaxone | 0
    initial treatment with clarithromycin | 0
    initial treatment with hydroxychloroquine | 0
    initial treatment with enoxaparin s.c. 40 mg once daily | 0
    progressed to hypoxaemic respiratory failure | 24
    trachea intubated | 24
    connected to ventilation | 24
    developed obstructive shock | 72
    echocardiography demonstrated severe right ventricular dysfunction | 72
    echocardiography demonstrated right atrial thrombus | 72
    received veno:arterial ECMO | 72
    received catheter-directed thrombolysis alteplase infusion | 72
    right ventricular function improved | 96
    right atrial thrombus disappeared | 96
    ECMO removed | 144
    CT pulmonary angiography confirmed pulmonary embolism | 144
    chest CT indicated COVID-19 pneumonia | 144
    weaned from ventilation | 192
    discharged from the hospital | 0
    received vitamin K antagonist | 0
    overlapping period with LMWH | 0
    follow-up echocardiography after 30 days showed mild pulmonary hypertension | 720
    follow-up echocardiography after 30 days showed normal right ventricle | 720
    rehabilitation programme as inpatient | 0
    good physical improvement | 0
    no neurological sequelae | 0
    no bleeding complications | 0
    <|eot_id|>