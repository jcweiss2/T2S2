40-day-old | 0
male | 0
neonate | 0
admitted to the hospital | 0
tricuspid valve mass | 0
neonatal seizures | -480
necrotizing enterocolitis | -480
blood cultures done | -480
anti-convulsants | -480
intravenous antibiotics | -480
piperacillin tazobactam combination | -480
amikacin | -480
peripheral venous access | -480
echocardiography done | -480
tricuspid mass | -480
referred to our centre | -20
not febrile | 0
deeply icteric | 0
no focal neurologic deficits | 0
no clinical heart failure | 0
clinical cardiovascular examination normal | 0
cephalhematoma | 0
computed tomography brain scan | 0
small petechial hemorrhages | 0
no space occupying lesions | 0
echocardiography showed vegetation | 0
vegetation attached to the tricuspid valve | 0
Doppler examination showed mean tricuspid inflow gradient | 0
blood cultures collected | 0
fungal cultures grew white yeast-like colonies | 24
organism identified as K. ohmeri | 24
Gram staining showed oval budding yeast cells | 24
antifungal susceptibility test | 24
MIC of anti-fungal agents | 24
amphotericin B started | 24
intravenous amphotericin B | 24
packed cell transfusion | 24
planned for surgical removal of the mass | 24
hemodynamic compromise | 48
fungal septicemia | 48
could not be resuscitated | 48
died | 48