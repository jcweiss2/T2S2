seven years old | 0 | 0 | Factual
male | 0 | 0 | Factual
admitted to the hospital | 0 | 0 | Factual
pre-B-ALL | -672 | 0 | Factual
first relapse of pre-B-ALL | -168 | -168 | Factual
allogeneic HSCT | -168 | -168 | Factual
hemoglobin 8.5 g/dl | 0 | 0 | Factual
thrombocytes 13,000/μl | 0 | 0 | Factual
WBC 940/μl | 0 | 0 | Factual
neutrophils 50/μl | 0 | 0 | Factual
CRP 6.83 mg/dl | 0 | 0 | Factual
ferritin 182 μg/dl | 0 | 0 | Factual
cachexia | 0 | 0 | Factual
dry skin | 0 | 0 | Factual
pallor | 0 | 0 | Factual
multiple hematomas | 0 | 0 | Factual
hepatosplenomegaly | 0 | 0 | Factual
antibiotic, antiviral, and antifungal chemoprophylaxis | 0 | 168 | Factual
ceftriaxone | 0 | 168 | Factual
teicoplanin | 0 | 168 | Factual
acyclovir | 0 | 168 | Factual
caspofungin | 0 | 168 | Factual
pain in the left flank | 0 | 120 | Factual
morphine | 0 | 120 | Factual
somnolent and sleepy | 120 | 120 | Factual
cerebral side effect of blinatumomab | 120 | 120 | Possible
cerebral CT scan | 120 | 120 | Factual
MRI scan | 120 | 120 | Factual
multiple cerebral hemorrhages | 120 | 120 | Factual
cardio-respiratory decompensation | 120 | 120 | Factual
mechanical ventilation | 120 | 168 | Factual
catecholamine therapy | 120 | 168 | Factual
blinatumomab treatment stopped | 120 | 120 | Factual
hemoglobin 6.7 g/dl | 120 | 120 | Factual
thrombocytes 49,000/μl | 120 | 120 | Factual
WBC 120/μl | 120 | 120 | Factual
neutrophils 20/μl | 120 | 120 | Factual
CRP 23.13 mg/dl | 120 | 120 | Factual
ferritin 1439 μg/dl | 120 | 120 | Factual
multiple thrombi in the left and right ventricle | 120 | 120 | Factual
thromboembolic events | 120 | 120 | Factual
endocarditis | 120 | 120 | Possible
septic embolisms | 120 | 120 | Possible
meropenem | 120 | 168 | Factual
gentamicin | 120 | 168 | Factual
CT scans of the thorax, abdomen and pelvis | 132 | 132 | Factual
multiple, systemic thromboembolic lesions | 132 | 132 | Factual
ischemia | 132 | 132 | Factual
bleeding | 132 | 132 | Factual
infarction | 132 | 132 | Factual
bone marrow aspiration | 132 | 132 | Factual
bone marrow aplasia | 132 | 132 | Factual
lymphatic blasts | 132 | 132 | Factual
cerebral pressure rising | 132 | 168 | Factual
cerebral herniation | 168 | 168 | Factual
death | 168 | 168 | Factual
invasive mycosis of R. pusillus | 0 | 168 | Factual
autopsy | 168 | 168 | Factual
R. pusillus identified via PCR-based methods | 168 | 168 | Factual
disseminated infection | 0 | 168 | Factual
mucormycosis | 0 | 168 | Factual