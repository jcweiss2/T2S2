76 years old | 0
man | 0
psoriasis | 0
chronic kidney disease stage 4 | 0
creatinine clearance of 29 ml/min/1.73 m2 | 0
essential hypertension | 0
amlodipine | 0
atenolol | 0
admitted to the Emergency Department | 0
lowered level of awareness | 0
sustained bradycardia | 0
denied syncope | 0
denied angina | 0
denied palpitation | 0
heart rate of 26 beats per minute | 0
blood pressure of 80/40 mmHg | 0
mean arterial pressure of 53 mmHg | 0
body temperature of 35.6°C | 0
respiratory rate of 18 breaths per minute | 0
95% peripheral oxygen saturation | 0
physical examination unremarkable | 0
white blood cell count of 5.450 cells/μL | 0
creatinine level of 3.7 mg/dL | 0
serum potassium level of 7.3 mg/dL | 0
TSH of 4.92 μUI/mL | 0
C-reactive protein of 48.9 mg/dL | 0
chest X-ray normal | 0
transthoracic echocardiography normal systolic function | 0
transthoracic echocardiography normal diastolic function | 0
transthoracic echocardiography no remarkable changes with the heart valves | 0
left ventricular dimension 46 mm | 0
interventricular septum 9 mm | 0
posterior wall 9 mm | 0
ejection fraction 64% | 0
sinus bradycardia | 0
junctional escape rhythm | 0
BRASH syndrome considered | 0
intravenous bolus of sodium chloride 0.9% | 0
atropine | 0
glucagon | 0
calcium gluconate | 0
hydrocortisone | 0
sodium bicarbonate | 0
dextrose 20% with regular insulin | 0
previous medications suspended | 0
blood pressure maintained at <65 mmHg | 0
continuous infusion of epinephrine | 0
temporary transvenous pacemaker placed | 0
hyperkalemia corrected | 24
creatinine levels returned to baseline | 24
epinephrine infusion suspended | 96
temporary pacemaker removed | 120
sinus rhythm with heart rate of 60–70 bpm | 120
discharged | 192
ECG normal sinus rhythm | 192
serum creatinine 2.36 mg/dL | 192
potassium 4.9 mg/dL | 192
beta-blockers avoided | 192
BRASH syndrome diagnosed | 0
bradycardia | 0
renal failure | 0
AV nodal-blocking agents | 0
shock | 0
hyperkalemia | 0
hypovolemia | 0
transvenous pacing | 0
hemodialysis | 0
sepsis | 0
acute heart disease | 0
chronic renal failure | 0
beta-blocker use | 0
hyperkalemia component | 0
ECG findings bradycardia | 0
hemodynamic support | 0
correction of hyperkalemia | 24
beta-blocker withdrawal | 0
renal replacement therapy | 0
temporary transvenous pacemaker | 0
epinephrine continuous infusion | 0
multiple-organ failure | 0
death | 0
