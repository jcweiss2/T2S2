58 years old | 0
female | 0
admitted to the hospital | 0
fever | -240
fatigue | -240
generalized body aches | -240
diarrhea | -72
chest tightness | -72
shortness of breath | -72
leukopenia | -240
thrombocytopenia | -240
antibiotics | -240
antipyretics | -240
temperature 36.5 ℃ | 0
heart rate 117/min | 0
respiratory rate 45/min | 0
blood pressure 170/100 mmHg | 0
conscious state | 0
crackles in both lungs | 0
scattered skin petechiae | 0
swollen lymph node | 0
leukopenia | 0
thrombocytopenia | 0
elevated liver enzymes | 0
elevated muscle enzymes | 0
inflammatory indicators | 0
urine occult blood | 0
urine protein | 0
pulmonary infection | 0
sepsis | 0
empiric antibiotic treatment | 0
biapenem | 0
voriconazole | 0
mental confusion | 24
endotracheal intubation | 24
mechanical ventilation | 24
serological tests | 24
serum galactomannan | 24
1,3-β-d-glucan | 24
mNGS | 24
Aspergillus fumigatus | 24
Aspergillus flavus | 24
Aspergillus terreus | 24
SFTSV | 24
ribavirin | 24
transfusion of plasma | 24
transfusion of platelet | 48
acute renal failure | 48
heart failure | 48
CRRT | 48
metaraminol | 48
fever | 168
leukocytosis | 168
procalcitonin | 168
Acinetobacter baumannii | 168
tigecycline | 168
pulmonary function improved | 216
radiological findings improved | 216
limb twitching | 408
thrombocytopenia | 408
anemia | 408
elevated creatine kinase | 408
prolonged activated partial thromboplastin time | 408
uncontrolled white mold | 408
repeat mNGS | 408
A. fumigatus | 408
discharged home | 432
died | 438