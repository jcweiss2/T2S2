32 years old | 0
male | 0
Caucasian | 0
admitted to the hospital | 0
epigastric pain | -48
ruptured appendicitis | -48
laparoscopic appendectomy | -48
fevers | -168
abdominal pain | -168
severe right upper quadrant epigastric pain | -168
septic shock | -168
temperature 103°F | -168
pulse 108 beats/minute | -168
mean arterial pressure of 47 mmHg | -168
fluid resuscitation | -168
vasopressors | -168
vancomycin | -168
piperacillin/tazobactam | -168
elevated white blood cell count | -168
absolute neutrophil count of 12,400 cells/mm^3 | -168
splenomegaly | -168
acute thrombosis of the proximal main portal vein | -168
Fusobacterium necrophorum | -168
metronidazole | -144
anticoagulation with intravenous heparin | -144
abdominal pain persisted | -120
thrombus continued to progress | -120
venography | -120
cavernous transformation of the portal vein | -120
transhepatic endovascular thrombolysis | -96
tissue plasminogen activator (tPA) | -96
recanalizing the porto-mesenteric veins | -96
discharged home | 168
warfarin | 168
oral clindamycin | 168
complete symptom relief | 336