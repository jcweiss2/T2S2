21 years old | 0
male | 0
obese | 0
admitted to the hospital | 0
cough | -72
fever | -72
shortness of breath | -72
pleuritic chest pain | -72
light-headedness | -72
near syncope | -72
dyspnoea | -72
COVID-19 | 0
sub-massive pulmonary embolism | 0
unfractionated heparin | 0
hypotensive | 12
massive pulmonary embolism | 12
catheter-directed thrombolysis | 12
improved clinically | 24
discharge planned | 24
acute respiratory failure | 96
hypotension | 96
intubated | 96
cardiac arrest | 96
return of spontaneous circulation | 96
vasopressors | 96
extracorporeal membrane oxygenation | 96
recurrent massive pulmonary embolism | 96
repeat catheter-directed thrombolysis | 96
ventilation parameters improved | 144
vasopressors discontinued | 144
weaning of ECMO | 144
deep venous thrombus | 144
inferior vena cava filter | 144
low-molecular-weight heparin | 144
septic shock | 240
treated with broad spectrum antibiotics | 240
right thigh haematoma | 240
compartment syndrome | 240
surgical debridement | 240
transitioned to rivaroxaban | 240
discharged to an acute rehabilitation facility | 1248
returned home | 1608
performing activities of daily living independently | 1608
anticoagulated on rivaroxaban | 1608
no major adverse events | 1608