12 years old | 0  
    female | 0  
    behavioural change | -144  
    fever | -144  
    headache | -144  
    conversation with self | -168  
    crying or laughing without reason | -168  
    altered consciousness | -168  
    abnormal hand movements | -168  
    inability to write letters | -168  
    sleep disturbance | -168  
    aggressive behaviour | -96  
    incomprehensive language | -96  
    visual hallucinations | -96  
    intermittent screaming | -96  
    high-grade fever | -96  
    admitted to Hua Hin Hospital | -96  
    ceftriaxone | -96  
    acyclovir | -96  
    azithromycin | -96  
    oseltamivir | -96  
    referred to King Chulalongkorn Memorial Hospital | 0  
    low-grade fever | 0  
    confusion | 0  
    disorientation | 0  
    oromotor dyskinesia | 0  
    choreoathetosis | 0  
    positive NMDAR autoantibodies | 0  
    generalized slow waves on EEG | 0  
    delta brush pattern on EEG | 0  
    seizure | 0  
    status epilepticus | 0  
    pulse methylprednisolone | 0  
    intravenous immunoglobulin | 0  
    prednisolone | 0  
    upper gastrointestinal bleeding | 1008  
    bilious vomiting | 1008  
    abdominal distension | 1008  
    watery diarrhoea | 1008  
    stool mixed with blood | 1008  
    Pseudomonas aeruginosa in stool | 1008  
    CMV PCR positive | 1008  
    CMV esophago$enterocolitis | 1008  
    ganciclovir | 1008  
    repeated pulse methylprednisolone | 1008  
    diarrhoea subsided | 1512  
    vomiting subsided | 1512  
    normal mucosa on endoscopy | 1512  
    cyclophosphamide | 1512  
    neurological improvement | 1512  
    discharged | 1512  
