40 years old | 0
male | 0
presented with a 4-day history of fever | -96
nausea | -96
vomiting | -96
enlarging non-tender left neck swelling | -96
hypotensive | 0
febrile | 0
confused | 0
unilateral anterior cervical triangle swelling | 0
erythematous rash on the left side of his neck | 0
erythematous rash on the anterior chest wall | 0
sinus rhythm | 0
left anterior fascicular block | 0
intravenous fluid resuscitation | 0
broad-spectrum antibiotics | 0
elevated CRP | 0
acute inflammatory process of the left submandibular space | 0
unilateral enlarged lymph nodes | 0
necrotizing lymphadenopathy | 0
clinical deterioration | 0
admission to ICU | 0
septic shock | 0
normal haemoglobin | 0
elevated neutrophils | 0
elevated inflammatory markers | 0
lymphopoenia | 0
thrombocytopoenia | 0
hyponatraemia | 0
hepatitis | 0
hypoalbuminaemia | 0
coagulopathy | 0
myocarditis | 0
negative viral and bacterial investigations | 0
negative vasculitis screen | 0
normal left ventricular function | 0
moderate central mitral regurgitation | 0
ongoing broad-spectrum antibiotics | 0
critically unwell | 0
ultrasound-guided biopsy of left anterior cervical lymph node on Day 3 | 72
suppurative necrotizing lymphadenitis | 72
new erythema of the oral mucosa on Day 4 | 96
fissured lips on Day 4 | 96
strawberry tongue on Day 4 | 96
bilateral conjunctival injection on Day 4 | 96
persistent fever | 96
diagnosis of classic Kawasaki disease | 96
treatment with IVIG | 96
high-dose aspirin | 96
clinical improvement within 2 days | 168
acute transient left upper limb weakness on Day 10 | 240
CT angiogram | 240
MRI | 240
excluded vertebral artery dissection | 240
excluded stroke | 240
CTCA at 3 months | 2160
two sequential aneurysms in RCA | 2160
aneurysm in LAD | 2160
no thrombus | 2160
no mural thickening | 2160
no coronary plaque | 2160
no perivascular fatty changes | 2160
cardiac MRI showed normal left ventricular volumes | 2160
preserved function | 2160
mid-wall fibrosis | 2160
follow-up CTCA at 12 months | 8760
resolution of LAD aneurysm | 8760
improvement of RCA aneurysms | 8760
