67 years old | 0
male | 0
admitted to the hospital | 0
dyspnea | 0
chest pain | 0
tachycardic | 0
tachypneic | 0
hypotensive | 0
elevated WBC count | 0
lactic acid elevated | 0
liver enzymes elevated | 0
electrocardiography showed sinus tachycardia with low voltage | 0
intubated | 0
pericardiocentesis | 0
removal of 800 mL of cloudy, milky fluid | 0
admitted to the ICU | 0
provisional diagnosis of rheumatoid pericardial effusion | 0
cardiac tamponade | 0
septic shock | 0
aggressively resuscitated | 0
pressor support | 0
broad-spectrum antibiotics | 0
blood and urine cultures were negative | 0
indium scan | 0
WBC accumulation within the upper abdomen | 0
discharged to a skilled nursing facility | 24
returned to the ED | 168
recurrent shortness of breath | 168
moderate pericardial effusion | 168
pericardial window | 168
generalized abdominal and back pain | 168
recurrent leukocytosis | 168
elevated lipase | 168
CT demonstrated a gas-containing fluid collection | 168
surgical exploration of the subxiphoid window | 168
pancreaticopericardial fistula | 168
infected pericardial window | 168
irrigate the pericardial space | 168
place a drain | 168
increasingly jaundiced | 192
wound infection | 192
enzymatic breakdown | 192
wound vacuum | 192
somatostatin | 192
EGD | 192
ERCP | 192
organized necrosis | 192
communication to the lumen | 192
side branch disruption | 192
pancreatic duct stent | 192
hypotensive | 216
unable to maintain adequate perfusion | 216
emergent family meeting | 216
limit treatment to comfort measures | 216
expired | 216
rheumatoid arthritis | -10080
tocilizumab | -10080 
severe rheumatoid arthritis | -10080