37 years old | 0
male | 0
healthcare worker | 0
close contact with COVID-19 patient | -120
high-grade fever | -96
myalgia | -96
dry cough | -96
tested positive for COVID-19 | -72
self-isolate at home | -72
worsening shortness of breath | -48
admitted to hospital | 0
bibasal crackles | 0
gallop rhythm of the heart | 0
resting tachycardia | 0
no signs of pedal oedema | 0
lymphopaenia | 0
raised C reactive protein | 0
lactate dehydrogenase | 0
brain natriuretic peptide | 0
mildly deranged liver function tests | 0
cardiac troponins negative | 0
ECG showed sinus tachycardia | 0
chest X-ray showed minimal bibasal infiltrates | 0
transthoracic echocardiogram | 0
eyeball ejection fraction estimate of 10%–15% | 0
dilated left ventricle | 0
left ventricular dimensions calculated | 0
serial cardiac troponins | 0
serial ECGs | 0
serial TTE | 0
gradual improvement in ejection fraction | 168
shortness of breath improved | 168
cardiac MRI | 504
moderate LV impairment | 504
no obvious evidence for myocardial fibrosis | 504
high-grade temperature spikes | 0
CRP <100 mg/L | 0
ceftriaxone prescribed | 0
blood and urine cultures negative | 0
CRP started creeping up | 72
ceftriaxone changed to piperacillin/tazobactam and vancomycin | 72
renal functions started deteriorating | 120
vancomycin stopped | 120
renal replacement therapy | 168
renal biopsy | 168
acute tubular injury | 168
granular casts | 168
localised inflammation around injured tubules | 168
intermittent haemodialysis | 168
significant improvement prior to discharge | 336
ejection fraction increased to 25%–30% | 336
renal function improving | 336
discharged | 336
follow-up cardiac MRI | 744
ejection fraction of 46% | 744
moderate LV impairment | 744
renal function within normal range | 744