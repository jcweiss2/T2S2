30 years old | 0
male | 0
no past medical history | 0
admitted to cardiac intensive care unit | 0
second dose of mRNA SARS-CoV-2 vaccine | -40
fever | -39
pleuritic chest pain | -39
reduction of symptoms | -35
presyncope | -10
hospital admission | -10
diagnosis of acute pericarditis | -10
cardiac tamponade | -10
pericardiocentesis | -10
non-steroid anti-inflammatory drugs | -10
colchicine | -10
symptom remission | -3
inflammatory markers downward trend | -3
discharge | -3
relapse of pleuritic chest pain | 8
elevated inflammatory markers | 8
moderate pericardial effusion | 8
admitted to Cardiology ward | 8
worsening pericardial effusion | 10
mild signs of impaired ventricular filling | 10
C-reactive protein 306 mg/L | 10
anakinra started | 10
no chest pain | 11
C-reactive protein 287 mg/L | 11
no chest pain | 12
C-reactive protein 179 mg/L | 12
complete reabsorption of pericardial effusion | 13
C-reactive protein 104 mg/L | 13
C-reactive protein 34 mg/L | 15
discharge | 16
asymptomatic | 16
good clinical conditions | 16
anakinra 100 mg/day | 16
ibuprofen 600 mg t.i.d. | 16
colchicine 0.5 mg b.i.d. | 16
proton pump inhibitor | 16
follow-up visit | 28
asymptomatic | 28
telephonic contact | 60
asymptomatic | 60