39 years old | 0
female | 0
height 155 cm | 0
weight 44.5 kg | 0
mild dyspnea | 0
adenoid cystic carcinoma in the carina | 0
carinal resection and reconstruction | 0
left mainstem bronchus almost totally obstructed | 0
mass extended to the carina and right mainstem bronchus | 0
internal diameter of the RMB 11 mm | 0
length of the RMB 12 mm | 0
length of the distal LMB not involved by the mass 20 mm | 0
no underlying diseases | 0
preoperative examinations normal findings | 0
moderate obstructive pattern of the pulmonary function test | 0
forced expiratory volume in one second 1.88 liter | 0
forced vital capacity 2.81 liter | 0
ratio 67% | 0
general anesthesia induced | 0
target-controlled infusion of propofol | 0
target-controlled infusion of remifentanil | 0
rocuronium 40 mg | 0
tracheal intubation | 0
right-sided double-lumen tube | 0
patient moved to the right lateral position | 0
left bronchi and vasculature dissected | 0
thoracoscopic surgery under right OLV | 0
arterial oxygen tension 462 mmHg | -20
inspired oxygen fraction 1.0 | -20
right-sided double-lumen tube replaced | 0
single-lumen endotracheal tube | 0
bronchial blocker | 0
patient moved to the left lateral position | 0
right thoracotomy | 0
peak airway pressure 28 cmH2O | 0
tidal volume 300 ml | 0
arterial oxygen tension 110 mmHg | 20
inspired oxygen fraction 1.0 | 20
carinal resection | 0
LMB resected | 0
sterile reinforced endotracheal tube | 0
left OLV | 0
airway pressure 35 cmH2O | 0
oxygen saturation 70% | 0
RMB resected | 0
additional sterile endotracheal tube | 0
differential bilateral lung ventilation | 0
oxygen saturation 100% | 2
carina removed | 0
RMB anastomosed with the resected trachea | 0
no air leak | 0
LMB implanted to neither the trachea nor the right bronchus | 0
left lung removed | 0
left endobronchial tube removed | 0
non-dependent right lung ventilated | 0
low tidal volume 200-250 ml | 0
airway pressure lower than 20 cmH2O | 0
oxygen saturation below 80% | 0
tube reinserted into the LMB | 0
two-lung ventilation | 0
right OLV reattempted | 0
oxygen saturation below 90% | 3
left pulmonary artery clamped | 0
right OLV attempted | 0
oxygen saturation 100% | 5
left main pulmonary artery ligated | 0
left endobronchial tube removed | 0
right thoracotomy closed | 0
patient moved to the right lateral position | 0
left thoracotomy | 0
left pulmonary artery and veins resected | 0
left pneumonectomy | 0
patient shifted to the supine position | 0
chin tightly sutured to the chest | 0
tracheal extubation | 0
patient transferred to the intensive care unit | 0
discharged on the 13th postoperative day | 312