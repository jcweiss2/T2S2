28 years old | 0
male | 0
admitted to the hospital (burn intensive care unit) | 0
mixed partial-thickness burns | 0
full-thickness burns | 0
53% total body surface area burns | 0
burns to face | 0
burns to chest | 0
burns to bilateral upper extremities | 0
burns to bilateral lower extremities | 0
burns to abdomen | 0
intubated | 0
minimal ventilatory support | 0
oxygen saturation (Spo2) of 100% | 0
arterial partial pressure of oxygen (Pao2) of 326 mm Hg | 0
crystalloid fluid resuscitation | 0
titrated fluid resuscitation | 0
urine output monitoring | 0
acutely worsening hypoxemia | -72
escalation of inspired oxygen fraction (Fio2) | -72
high positive end-expiratory pressure | -72
sedation | -72
neuromuscular blockade | -72
respiratory status deterioration | -72
Pao2/Fio2 of 50 mm Hg | -72
chest radiograph on hospital day 3 | -72
bilateral pulmonary infiltrates | -72
ARDS | -72
emergent VV=ECMO initiation | -72
19-French reinfusion cannula placement | -72
23-French drainage cannula placement | -72
ECMO flows of 4.7 to 5.0 L/min | -72
transient Spo2 improvement >90% | -72
oxygenation status worsening | -24
Pao2/Fio2 of 43 mm Hg | -24
echocardiogram | -24
elevated cardiac output (10-11 L/min) | -24
ECMO flow limitation to 5 L/min | -24
suction events | -24
ECMO flow/native CO ratio of 0.45-0.50 | -24
strategies to reduce CO | -24
decreasing body temperature | -24
beta-blockade initiation | -24
unsuccessful CO reduction | -24
reinfusion cannula repositioning | -24
bilateral femoral vein drainage cannulas in Y configuration | -24
20-French reinfusion cannula placement | -24
veno-VV-ECMO reconfigured | -24
ECMO flows increased to 6-6.5 L/min | -24
hypoxemia persistence | -24
Pao2/Fio2 of 48 mm Hg | -24
elevated lactate dehydrogenase (>1400 units/L) | -24
multiple ECMO oxygenator exchanges | -24
postoxygenator Pao2 100-200 mm Hg | -24
second ECMO circuit insertion | 0
parallel VV-ECMO circuits | 0
combined flow of 6 L/min | 0
flow synchronization | 0
postoxygenator Pao2 >350 mm Hg | 0
Spo2 >90% | 0
lactate dehydrogenase decrease (<600 units/L) | 0
respiratory status improvement | 96
Pao2/Fio2 of 430 mm Hg | 96
heavy diuresis | 96
pulmonary hygiene | 96
ventilator settings weaned to Fio2 40% | 96
parallel VV-ECMO weaning | 96
one system weaned down | 96
ECMO decannulation | 240
sepsis | 240
pneumonia | 240
bacteremia | 240
fungemia | 240
gastrointestinal bleeding | 240
multiple debridements | 240
skin grafts | 240
discharged on room air | 2160
