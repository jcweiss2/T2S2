67 years old | 0
male | 0
admitted to the hospital | 0
untreated hypertension | 0
diabetes | 0
acutely increasing chest pain | -12
back pain | -12
ST segment elevation in V1-6 | 0
wall motion abnormality in the anterior region | 0
anterior acute STEMI diagnosis | 0
maximum creatinine kinase level 5021 U/L | 0
maximum CK-MB level 535 U/L | 0
coronary angiography revealed total occlusion at the middle section of the left anterior descending artery | 0
percutaneous coronary intervention performed | 0
chest pain occurred on a previous day | -36
CK level already high at admission | 0
acute strong right subcostal pain 5 hours after PCI | 5
acute strong epigastric pain 5 hours after PCI | 5
abdominal computed tomography performed | 5
acute cholecystitis suspected | 5
gallstones detected | 5
liver enzyme level did not increase | 5
treated conservatively for biliary colic | 5
no symptoms of left heart failure | 0
no dyspnea during exertion | 0
no orthopnea | 0
symptoms of right heart failure | 0
fatigue | 0
loss of appetite | 0
myocardial enzyme level decreased after PCI | 0
no heart murmur heard | 0
no evidence of new ECG abnormalities | 0
daily TTE did not demonstrate new signs of decreased systolic function | 0
daily TTE did not demonstrate new signs of myocardial ischemia | 0
daily TTE did not demonstrate new signs of mechanical complications | 0
stronger right subcostal pain on 5th day | 120
stronger epigastric pain on 5th day | 120
positive Murphy sign | 120
no heart murmur | 120
C-reactive protein increase to 10.82 mg/dL | 120
new CT revealed edematous gallbladder | 120
white blood cell count increased to 12600/µL | 120
aspartate aminotransferase 57 U/L | 120
alanine aminotransferase 45 U/L | 120
gamma-glutamyl transpeptidase 77 U/L | 120
gallstones vanished | 120
abdominal symptoms strongly suspicious of acute cholecystitis | 120
laparoscopic cholecystectomy performed | 120
chronic cholecystitis identified by pathological examination | 120
postoperative exacerbated pain | 120
admission to ICU due to restlessness | 144
tachypnea | 144
shock | 144
no new abnormality on TTE | 144
no new abnormality on ECG | 144
septic shock management | 144
broad-spectrum antibiotics | 144
tracheal intubation | 144
invasive ventilation | 144
continuous renal replacement therapy | 144
norepinephrine administration | 144
dobutamine administration | 144
epinephrine administration | 144
hemodynamic state deteriorated | 144
4 times TTE indicated no abnormalities after ICU admission | 144
5th TTE revealed left-to-right shunt through ventricular septum | 154
VSR suspected | 154
intra-aortic balloon pumping | 154
venous-artery extracorporeal membrane oxygenation | 154
emergency patch closure of VSR performed | 154
perforation at apical septal region confirmed by TEE | 154
perforation confirmed by surgeons’ inspection | 154
right subcostal pain diminished | 154
hemodynamics improved | 154
left ICU on 21st day | 504
transferred on 74th day | 1776
