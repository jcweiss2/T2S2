60 years old | 0
male | 0
hypertension | 0
unspecified left ventricular dysfunction | 0
chest pain | -285
beta-blockers | 0
sartanic | 0
tiazidic diuretic | 0
called emergency department | -15.5
awake | -15.5
hypotensive | -15.5
symptomatic | -15.5
ECG signs of extensive antero-lateral AMI | -15.5
morphine | -15.5
apirine | -15.5
dopamine infusion | -15.5
transferred to peripheral hospital | -15.5
angiographic study | -13.5
severe cardiogenic shock | -13.5
unresponsive to catecholamine | -13.5
IABP support | -13.5
distal occlusion of left main coronary artery | -13.5
angioplasty | -13.5
positioned bare metal stent | -13.5
heparin bolus 7500 IU | -13.5
continuous infusion of reopro | -13.5
good revascularization | -13.5
TIMI score 1 | -13.5
severe hypotension | -13.5
high-dose norepinephrine | -13.5
bradi-asystolic cardiac arrest | -12.5
advanced life support algorithms | -12.5
tracheal intubation | -12.5
transvenous pacing | -12.5
cardiogenic shock refractory | -12.5
high amines dosage | -12.5
mechanical ventilation | -12.5
systolic blood pressure 90 mmHg | -12.5
heart rate 100 beats per minute | -12.5
anuria | -12.5
paO2 53 mmHg | -12.5
paCO2 60 mmHg | -12.5
pH 7.04 | -12.5
lactates >6 mmol/L | -12.5
base excess -14 mmol/L | -12.5
echocardiography showed contractile reserve | -12.5
called ECMO team | -10
ECMO implantation | -8.75
percutaneous cannulation of right femoral artery | -8.75
percutaneous cannulation of left femoral vein | -8.75
ECMO circuit prepared | -8.75
connected to ECMO | -8
blood flow 3.5 L/min | -8
gas flow 3 L/min | -8
FiO2 0.6 | -8
hemodynamic stabilization | -8
reduction of amines | -8
recovery of diuresis | -8
normalization of blood gas parameters | -8
PaO2 457 mmHg | -8
PaCO2 29 mmHg | -8
pH 7.48 | -8
lactates 1,9 mmol/L | -8
BE -1,2 mmol/L | -8
reopro infusion interrupted | -8
transferred to San Gerardo Hospital | -7
sedated | 0
continuous perfusion of muscle relaxant | 0
therapeutic hypothermia | 0
hemodynamically stable | 0
arterial catheter | 0
central venous catheter | 0
pulmonary artery catheter | 0
arterial blood pressure 150/60 mmHg | 0
heart rate 80 beats | 0
sinus rhythm | 0
central venous pressure 12 mmHg | 0
wedge pressure 15 mmHg | 0
pulmonary artery pressure 29/18 mmHg | 0
cardiac output 2,5 L/min | 0
venous oxygen saturation 72% | 0
transesophageal echocardiography showed ejection fraction 10% | 0
dobutamine 5 mcg/kg/min | 0
intravenous heparin | 0
activated clotting time 180-200 seconds | 0
aspirin | 0
clopidrogel | 0
echocardiography showed akinesia | 24
daily evaluations of legs perfusion | 24
relative hypertension | 96
calcium-sensitizer infusion | 96
weaning from ECMO | 96
blood flow 2 L/min | 96
blood flow 1 L/min | 108
weaned from ECMO | 120
IABP | 120
dobutamine 10 mcg/kg/min | 120
cannulae removed | 120
hyperdynamic shock | 120
cardiac output 11 L/min | 120
blood pressure 80/40 mmHg | 120
norepinephrine | 120
treated as septic shock | 120
cultural examination | 120
empiric antibiotic therapy with meropenem | 120
removed IABP | 144
started nitrates | 144
echocardiography showed persisting akinesia | 144
ejection fraction 30% | 144
linezolid added | 168
fever | 168
elevation of leukocytes | 168
inflammation indexes | 168
bronchial bleeding | 168
deterioration of blood gas parameters | 168
high PEEP | 168
interruption of heparin | 168
interruption of clopidogrel | 168
Ecodoppler performed | 168
hypertensive crisis | 192
pulmonary oedema | 192
mechanical ventilation with PEEP 15cmH2O | 192
high FiO2 | 192
inhalatory nitric oxide | 192
negative water balance | 192
calcium-sensitizer infusion | 192
diastolic dysfunction | 192
ACE-inhibitor | 192
beta-blockers | 192
extubated | 264
digoxin introduced | 312
transferred back to original hospital | 480
awake | 480
no neurological deficits | 480
hemodynamically stable | 480
sinus rhythm | 480
ACE-inhibitor | 480
beta-blocker | 480
normal renal function | 480
normal blood gas analysis | 480
