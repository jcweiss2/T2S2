56 years old| 0
    male| 0
    chronic kidney disease| 0
    maintenance hemodialysis| 0
    septic shock| 0
    coagulopathy| 0
    dialysis catheter in right internal jugular vein| 0
    attempted cannulation of left internal jugular vein with triple-lumen central venous catheter| 0
    catheter malpositioned| 0
    transferred from dialysis unit to ICU| 0
    altered sensorium| 0
    hypotension| 0
    Glasgow coma scale score 7/15: E2, V2, M3| 0
    heart rate 112 beats/min| 0
    blood pressure 87/48 mmHg| 0
    axillary temperature 38.5℃| 0
    dialysis-related septic shock diagnosis| 0
    fluid resuscitation initiated| 0
    routine cultures initiated| 0
    empirical antibiotic therapy initiated| 0
    intubated electively| 0
    mechanical ventilation| 0
    leukocyte count 17 × 10^6/cm³| 0
    sodium 122 mEq/L| 0
    potassium 3.2 mEq/L| 0
    international normalized ratio 3.2| 0
    normal platelet count| 0
    vasopressor therapy considered| 0
    dialysis catheter in right IJV considered for vasopressors| 0
    nephrology team consultation| 0
    decision to place separate central venous catheter in left IJV| 0
    dialysis catheter considered sepsis source| 0
    ultrasound-guided insertion of catheter into left IJV| 0
    catheter insertion successful up to 12 cm mark| 0
    post-procedure chest X-ray showed catheter loop in left brachiocephalic vein| 0
    catheter tip in left subclavian vein| 0
    dialysis catheter in right IJV considered obstacle| 0
    dialysis catheter removed| 0
    new dialysis catheter placed in femoral vein| 0
    central line repositioned using guidewire| 0
    follow-up chest X-ray showed catheter in right subclavian vein| 0
    decision to withdraw catheter 1-2 cm| 0
    catheter tip placed at junction of great veins| 0
    discussion of central venous access urgency| 0
    consideration of using existing dialysis catheter| 0
    patient dependent on dialysis| 0
    dialysis catheter possibly infected| 0
    alternative sites considered: right/left subclavian, left IJV, femoral veins| 0
    subclavian approach avoided due to coagulation abnormalities| 0
    femoral vein CVP reliability controversy| 0
    femoral route complications considered| 0
    left IJV approach chosen| 0
    bilateral IJV cannulation risks considered| 0
    patient with possible decreased cerebral perfusion| 0
    left IJV cannulation with triple-lumen catheter opted| 0
    catheter misplacement discussed| 0
    left side catheterization challenges| 0
    ideal catheter tip position discussed| 0
    initial catheter loop formation explained| 0
    guidewire-assisted repositioning| 0
    dialysis catheter removal impact| 0
    catheter withdrawal to superior vena cava| 0
    ultrasound guidance benefits noted| 0
    catheter tip malposition inevitability acknowledged| 0
    best practice consideration: remove dialysis catheter first| 0
    inability to remove dialysis catheter initially| 0
    undetermined cause of catheter misplacement| 0
    fluoroscopy/venography considerations| 0
    patient condition restrictions| 0
    expedited radiographic confirmation recommended| 0
    serial X-rays emphasized| 0
    chest X-ray showing right IJV dialysis catheter and central venous catheter loop| 0
    chest X-ray after catheter repositioning| 0
    chest X-ray after catheter withdrawal| 0
    patient consented to case publication| 0
    <|eot_id|>
    56 years old|0
male|0
chronic kidney disease|0
maintenance hemodialysis|0
septic shock|0
coagulopathy|0
dialysis catheter in right internal jugular vein|0
attempted cannulation of left internal jugular vein with triple-lumen central venous catheter|0
catheter malpositioned|0
transferred from dialysis unit to ICU|0
altered sensorium|0
hypotension|0
Glasgow coma scale score 7/15: E2, V2, M3|0
heart rate 112 beats/min|0
blood pressure 87/48 mmHg|0
axillary temperature 38.5℃|0
dialysis-related septic shock diagnosis|0
fluid resuscitation initiated|0
routine cultures initiated|0
empirical antibiotic therapy initiated|0
intubated electively|0
mechanical ventilation|0
leukocyte count 17 × 10^6/cm³|0
sodium 122 mEq/L|0
potassium 3.2 mEq/L|0
international normalized ratio 3.2|0
normal platelet count|0
vasopressor therapy considered|0
dialysis catheter in right IJV considered for vasopressors|0
nephrology team consultation|0
decision to place separate central venous catheter in left IJV|0
dialysis catheter considered sepsis source|0
ultrasound-guided insertion of catheter into left IJV|0
catheter insertion successful up to 12 cm mark|0
post-procedure chest X-ray showed catheter loop in left brachiocephalic vein|0
catheter tip in left subclavian vein|0
dialysis catheter in right IJV considered obstacle|0
dialysis catheter removed|0
new dialysis catheter placed in femoral vein|0
central line repositioned using guidewire|0
follow-up chest X-ray showed catheter in right subclavian vein|0
decision to withdraw catheter 1-2 cm|0
catheter tip placed at junction of great veins|0
discussion of central venous access urgency|0
consideration of using existing dialysis catheter|0
patient dependent on dialysis|0
dialysis catheter possibly infected|0
alternative sites considered: right/left subclavian, left IJV, femoral veins|0
subclavian approach avoided due to coagulation abnormalities|0
femoral vein CVP reliability controversy|0
femoral route complications considered|0
left IJV approach chosen|0
bilateral IJV cannulation risks considered|0
patient with possible decreased cerebral perfusion|0
left IJV cannulation with triple-lumen catheter opted|0
catheter misplacement discussed|0
left side catheterization challenges|0
ideal catheter tip position discussed|0
initial catheter loop formation explained|0
guidewire-assisted repositioning|0
dialysis catheter removal impact|0
catheter withdrawal to superior vena cava|0
ultrasound guidance benefits noted|0
catheter tip malposition inevitability acknowledged|0
best practice consideration: remove dialysis catheter first|0
inability to remove dialysis catheter initially|0
undetermined cause of catheter misplacement|0
fluoroscopy/venography considerations|0
patient condition restrictions|0
expedited radiographic confirmation recommended|0
serial X-rays emphasized|0
chest X-ray showing right IJV dialysis catheter and central venous catheter loop|0
chest X-ray after catheter repositioning|0
chest X-ray after catheter withdrawal|0
patient consented to case publication|0

