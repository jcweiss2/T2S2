42 years old | 0
male | 0
admitted to the hospital | 0
fever | -72
cough | -72
dyspnoea | -72
headache | -72
diagnosed with COVID-19 | -72
RT-PCR was positive for SARS-CoV-2 | -72
trachea intubated | 24
connected to ventilation | 24
hypoxic respiratory failure | 24
echocardiography was normal | 0
obstructive shock | 72
severe right ventricular dysfunction | 72
right atrial thrombus | 72
veno-arterial extracorporeal membrane oxygenation (VA-ECMO) | 72
catheter-directed thrombolysis alteplase infusion | 72
right ventricular function improved | 96
right atrial thrombus disappeared | 96
ECMO was removed | 144
CT pulmonary angiography confirmed pulmonary embolism | 144
Chest CT indicated COVID-19 pneumonia | 144
weaned from ventilation | 192
discharged from the hospital | 720
moderate systolic hypertension | 0
heart rate of 94 b.p.m. | 0
respiratory rate of 30 breaths/min | 0
oxygen flow rate of 15 L/min | 0
O2 saturation of 94% | 0
no signs of left ventricular failure | 0
no leg oedema | 0
fine scattered crackles | 0
electrocardiogram (ECG) was normal | 0
echocardiogram on admission was normal | 0
Chest X-ray (CXR) showed bilateral peripheral pulmonary infiltrates | 0
white cell count of 19.5 × 109/L | 0
neutrophil count of 14.5 × 109/L | 0
lymphocyte count of 0.7 × 109/L | 0
platelet count of 360 × 109/L | 0
haematocrit of 24.6% | 0
ferritin level of 855 μg/L | 0
high-sensitivity C-reactive protein level of 112.0 mg/L | 0
D-dimer level of 4400 ng/mL | 0
fibrinogen level of 7.1 g/L | 0
prothrombin time of 17.0 s | 0
activated partial thromboplastin time (aPTT) of 43.7 s | 0
treated with ceftriaxone | 0
treated with clarithromycin | 0
treated with hydroxychloroquine | 0
treated with enoxaparin | 0
hypotension | 72
sinus tachycardia | 72
haemodynamically unstable | 72
ECG showed sinus tachycardia | 72
S1Q3T3 pattern | 72
acute T wave inversion | 72
point-of-care echocardiography evaluation showed a dilated and severely hypokinetic right ventricle | 72
mean derived pulmonary arterial pressure of 60 mmHg | 72
large mobile echogenic mass swirling around in the right atrium | 72
treated with high-dose norepinephrine | 72
treated with dobutamine | 72
treated with vasopressin | 72
started on VA-ECMO | 72
catheter-directed thrombolysis with alteplase infusion | 72
follow-up echocardiography showed a decrease in the right ventricular diameter | 96
improvement in systolic function | 96
decrease in pulmonary pressure | 96
disappearance of the clot | 96
VA-ECMO was removed | 144
CT scan of the chest revealed filling defects in the main left and right pulmonary arteries | 144
CT scan of the chest showed extensive multifocal areas of ground-glass opacities | 144
weaned from the ventilator | 192
started treatment with a vitamin K antagonist | 720
overlapping period with low molecular weight heparin (LMWH) | 720
discharged from the hospital with no symptoms | 720
follow-up echocardiography after 30 days showed mild pulmonary hypertension | 744
normal right ventricle | 744