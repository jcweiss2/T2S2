100-year-old | 0  
    male | 0  
    referred to emergency department | 0  
    anterior neck swelling | 0  
    dysphagia | 0  
    muffled voice | 0  
    presented to emergency department two weeks prior | -336  
    similar symptoms two weeks prior | -336  
    oral steroid | -336  
    presumed lymphadenitis | -336  
    symptoms did not abate with steroids | -336  
    unable to wear dentures for two weeks | -336  
    only could swallow liquids | 0  
    hyperlipidemia | 0  
    benign prostatic hyperplasia | 0  
    hypertension | 0  
    no history of alcohol use | 0  
    no history of tobacco use | 0  
    no history of illicit drug use | 0  
    physical exam | 0  
    no respiratory distress | 0  
    expressed discomfort secondary to pain | 0  
    heart rate 89 beats/min | 0  
    blood pressure 131/81 mmHg | 0  
    oxygen saturation 94% | 0  
    respiratory rate 18 breaths/min | 0  
    severely limited mouth-opening | 0  
    inter-incisor gap 1 cm | 0  
    unable to extend neck | 0  
    diffuse neck swelling | 0  
    neck pain | 0  
    white blood count 28,000/μL | 0  
    hemoglobin 12.1 g/dL | 0  
    platelet count 225,000/μL | 0  
    computerized tomography neck scan | 0  
    large peripherally enhanced loculated fluid collection | 0  
    surrounding soft tissue edema | 0  
    resilient mass effect | 0  
    narrowing of oropharynx | 0  
    no significant lymphadenopathy | 0  
    dental caries | 0  
    remaining three mandibular teeth | 0  
    lucency suggested dental abscess | 0  
    surgical drainage of abscess | 0  
    airway secured with awake fiberoptic intubation | 0  
    denitrogenated with 100% oxygen | 0  
    glycopyrrolate 0.2 mg | 0  
    nasal decongestant oxymetazoline 0.05% | 0  
    topical lidocaine | 0  
    positioned in seated position | 0  
    ketamine administered | 0  
    light sedation | 0  
    difficulty visualizing vocal cords | 0  
    endotracheal intubation successful | 0  
    placement of 7.5 mm cuffed endotracheal tube | 0  
    confirmation of endotracheal intubation | 0  
    fentanyl 50 mcg | 0  
    propofol 50 mg | 0  
    muscle relaxant not administered | 0  
    spontaneous breathing on ventilator | 0  
    sevoflurane | 0  
    dexamethasone 10 mg | 0  
    incision and drainage of abscess | 0  
    collection of cultures | 0  
    shifted to intensive care unit | 0  
    elective postoperative ventilation | 0  
    extubated successfully | 24  
    postoperative period | 24  
    surgical cultures revealed Streptococcus viridans | 24  
    surgical cultures revealed Streptococcus intermedius | 24  
    Ludwig’s angina | 0  
    airway soft tissue swelling | 0  
    edema | 0  
    deep neck space infection | 0  
    dental abscess | 0  
    anticipated difficult airway | 0  
    perioperative considerations | 0  
    multiple comorbidities | 0  
    poorer functional status | 0  
    frailty | 0  
    multi-disciplinary team approach | 0  
    life-threatening complications | 0  
    necrotizing fasciitis | 0  
    descending mediastinitis | 0  
    pleural effusion | 0  
    sepsis | 0  
    aspiration pneumonia | 0  
    risk of abscess rupture | 0  
    difficulty in ventilation | 0  
    difficulty in intubation | 0  
    anatomic changes in geriatric population | 0  
    decreased neck mobility | 0  
    impaired cough mechanism | 0  
    decreased ventilatory response | 0  
    decreased pulmonary reserve | 0  
    increased autonomic dysfunction | 0  
    impaired autoregulation | 0  
    malnutrition | 0  
    decreased compliance of submandibular space | 0  
    edentulousness | 0  
    airway collapse | 0  
    difficult seal with bag-valve-mask | 0  
    rapid diagnosis | 0  
    aggressive treatment | 0  
    appropriate antibiotic treatment | 0  
    perioperative neurocognitive dysfunction | 0  
    robust assessment of comorbidities | 0  
    risk stratification | 0  
    preoperative optimization | 0  
    rehabilitation | 0  
    discharge planning | 0  
    high-risk clinics | 0  
    comprehensive geriatric assessment | 0  
    vigilant management | 0  
    life-threatening emergency | 0  
    surgical airway | 0  
    less invasive methods | 0  
    risk-benefit ratio | 0  
    airway management plan | 0  
    decreased risk of airway collapse | 0  
    head in sniffing position | 0  
    maximal opening of pharyngeal airway | 0  
    accurate assessment of airway | 0  
    immediate confirmation of tube placement | 0  
    less sympathetic stimulation | 0  
    less risk for airway trauma | 0  
    polymicrobial infection | 0  
    Streptococcus species | 0  
    Peptostreptococcus species | 0  
    Bacteroides species | 0  
    anaerobes | 0  
    penicillin G | 0  
    metronidazole | 0  
    ampicillin-sulbactam | 0  
    clindamycin | 0  
    cefoxitin | 0  
    antibiotic regimen | 0  
    definitive management | 0  
    awake blind nasal intubation | 0  
    flexible fiberoptic nasal intubation | 0  
    oral intubation | 0  
    less invasive methods attempted | 0  
    surgical plan | 0  
    medical comorbidities | 0  
    clinical exam | 0  
    airway management plan discussed | 0  
    multi-disciplinary team discussion | 0  
    postoperative outcomes | 24  
    successful intubation | 0  
    successful surgical procedure | 0  
    successful postoperative ventilation | 24  
    successful extubation | 24  
    postoperative monitoring | 24  
    action plans implemented | 0  

