63 years old | 0
female | 0
admitted to the hospital | 0
history of transient ischemic attack | -672
history of reflux | -672
history of hypertension | -672
history of hyperlipidemia | -672
previous laparoscopic sleeve gastrectomy | -672
vitamin supplements | -672
weight loss | -672
weight gain | -168
worsening gastroesophageal reflux disease (GERD) symptoms | -24
esophagogastroduodenoscopy | -24
large hiatal hernia | -24
laparoscopic hand-assisted hiatal hernia repair | 0
conversion of sleeve gastrectomy to Roux-en-Y gastric bypass (RYGB) | 0
vast adhesive disease | 0
discharged home | 96
followed up at outpatient bariatric institute | 192
shortness of breath | 432
left lower leg pain | 432
swelling | 432
hypotensive | 432
unresponsive | 432
cardiopulmonary arrest | 432
cardiopulmonary resuscitation | 432
intubated | 432
admitted to ICU | 432
extremely acidotic | 432
acute hypoxic respiratory failure | 432
renal failure | 432
computed tomography (CT) imaging | 432
pulmonary embolism protocol | 432
enlarged left common iliac, external iliac, and common femoral veins | 432
edema of the left thigh | 432
therapeutic anticoagulation | 432
vascular surgery consultation | 432
substantial swelling | 432
purple discoloration | 432
cold to touch | 432
combined diagnostic laparoscopy and lower-extremity venogram | 432
diagnostic laparoscopy | 432
pink viable bowel | 432
no identified abnormalities | 432
venogram | 432
extensive, acute, nearly occlusive left iliac and femoral venous thrombosis | 432
clot retrieval system | 432
thrombectomy | 432
multisystem organ failure | 480
shock | 480
liver failure | 480
respiratory failure | 480
disseminated intravascular coagulation | 480
increasing vasopressor support | 480
significant acidosis | 480
continuous renal replacement therapy | 480
tense left lower extremity | 504
bullous formation of the skin | 504
mottled digits | 504
no identifiable pulses or Doppler signals | 504
compartment syndrome | 504
4-compartment calf fasciotomy | 504
viable muscle | 504
no abnormality | 504
fasciotomy | 504
copious brown fluid | 504
pale, unresponsive muscle | 504
tissue death | 504
cardio-pulmonary arrest | 528
resuscitation | 528
death | 528