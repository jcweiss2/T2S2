54 years old | 0
male | 0
insulin dependent diabetes mellitus | -672
hepatitis C chronic infection | -672
liver cirrhosis child B | -672
esophageal varices | -672
right sided facial weakness | 0
right sided headache | 0
blocked right nostril | 0
fever | -168
admitted to the hospital | 0
BP 140/70 mmHg | 0
Pulse of 92 beat per minute | 0
oxygen saturation on an ambient air of 99% | 0
Temperature of 38.2 Celsius | 0
conscious | 0
alert | 0
oriented | 0
no apparent distress | 0
swelling of the right side of the face | 0
right eye complete ptosis | 0
chemosis | 0
injection | 0
mid dilated fixed pupil | 0
right frozen globe | 0
multiple cranial nerves palsies | 0
II palsy on right side | 0
III palsy on right side | 0
IV palsy on right side | 0
V1 palsy on right side | 0
VI palsy on right side | 0
VII palsy on right side | 0
no other focal neurological deficits | 0
right central retinal artery occlusion | 0
edematous retina | 0
black discoloration in the roof of the nasal cavity | 0
pale mucosa | 0
high WBC count | 0
hyperglycemia | 0
abnormal kidney function | 0
pansinusitis | 0
IV fluids | 0
insulin | 0
IV liposomal amphotericin | 0
Linezolid | 0
ceftazidime | 0
right radical endoscopic sinus surgery | 24
wide debridement | 24
extubated | 24
stayed in the surgical intensive care | 24
CT head with Iodine based IV injection of medium contrast | 24
inflammatory changes of the optic nerve | 24
inflammatory changes of adjacent muscles | 24
bony defect in the right lamina papyracea | 24
nasal swab by microscopy returned positive for Mucor species | 24
histopathology confirmed the diagnosis of invasive mucormycosis | 96
afebrile | 96
blood sugar improved | 96
kidney function improved | 96
rose again | 96
serum creatinine 260 µmol/L | 96
amphotericin toxicity | 96
contrast induced nephropathy | 96
IV fluids support continued | 96
IV amphotericin continued | 96
decreased level of consciousness | 192
confusion | 192
drop of GCS to 9/15 | 192
stable vital signs | 192
management for presumed hepatic encephalopathy | 192
lactulose | 192
broad spectrum antibacterial agents | 192
monitoring of mental status | 192
level of consciousness didn’t improve | 192
brain MRI | 360
total occlusion of the right internal carotid artery | 360
right anterior and middle cerebral arteries causing edema effect | 360
compression of the right posterior cerebral artery | 360
secondary massive infarction | 360
whole right cerebral hemisphere | 360
upper brain stem | 360
left frontal and basal ganglia regions | 360
right cerebellar hemisphere | 360
evidence of hemorrhagic change | 360
secondary mass effect | 360
significant midline shift | 360
declared brain dead | 408
apnea test was positive | 408
thorough discussion with the family for withdraw of care | 408
family objected | 408
passed away | 504
refractory septic shock | 504