24 years old | 0
female | 0
right groin pain | -672
nightly pain | -168
sweating | -168
no prior history of hip pathology | 0
healthy | 0
contact sports | 0
no medications | 0
no intravenous drug use | 0
no smoking | 0
no immune suppression | 0
afebrile | 0
vital stability | 0
antalgic gait | 0
leg in slight flexion | 0
external rotation at rest | 0
internal rotation of hip tender | 0
restricted internal rotation of hip | 0
normal serum white cell count | 0
elevated C-reactive protein levels | 0
CT scan suggestive of pyomyositis | 0
no osseous destruction | 0
MRI revealed multiple abscesses | 0
small right hip joint effusion | 0
synovial enhancement | 0
antibiotic therapy withheld | 0
general anesthesia | 0
lateral decubitus position | 0
perineal post placement | 0
genitalia padded | 0
hip distracted | 0
surgical area prepped and draped | 0
anterolateral portal placement | 0
distal midanterior portal placement | 0
interportal capsulotomy | 0
hip distended with saline | 0
diagnostic arthroscopy | 0
purulence | 0
inflamed synovia | 0
synovial samples collected | 0
synovectomy | 0
psoas muscle release | 0
debridement of obturator externus | 0
obturator membrane pierced | 0
hole enlarged | 0
30-degree scope used | 0
intrapelvic abscess decompressed | 0
obturator internus debrided | 0
copious irrigation | 0
capsulotomy left open | 0
toe-touch weight bearing | 24
abduction brace | 24
afebrile postoperatively | 24
stable postoperatively | 24
CRP level 188 | 24
intraoperative cultures negative | 24
cefazolin IV | 24
discharged | 96
surgical pain at 3 weeks | 504
brace discontinued | 504
physiotherapy referral | 504
nontender at 6 weeks | 1008
hip flexor weakness | 1008
hip range of motion improved | 1008
CRP normalized | 1008
asymptomatic at 6 months | 4320
hip flexor strength regained | 4320
internal rotation improved | 4320
CRP normal | 4320
recurrence of abscess | 7200
right buttock pain | 7200
antalgic gait recurrence | 7200
limited hip range of motion | 7200
CRP level 70 | 7200
MRI showed abscess recurrence | 7200
open irrigation and debridement | 7200
