70 years old | 0
male | 0
Caucasian | 0
BMI 31.14 | 0
smoker | 0
hypertensive | 0
admitted to the hospital | 0
endovascular-aortic aneurysm repair | -2160
nephrectomy for kidney cancer | -2160
incisional hernia | -2160
laparoscopic treatment | -2160
multilayered mesh | -2160
follow-up | -720
CT scan | -720
endoleak from the aortic aneurysm | -720
recurrent incisional hernia | -720
aorto-bi-iliac bypass | -720
abdominal wall sublay prosthetic repair | -720
composite mesh | -720
partial resection of ileum | -720
removal of previously positioned mesh | -720
discharged | -672
US scan | -672
large periprosthetic haematoma | -672
percutaneous treatment with two drains | -672
drains removed | -665
fever | -662
leakage of enteric material | -662
CT scan | -662
diploid-pubic fluid collection | -662
jejunal fistula | -662
conservative management | -662
US guided positioning of two drains | -662
evacuation of 1800 cc of enteric material | -662
nasogastric tube | -662
total parenteral nutrition | -662
intravenous octreotide | -662
antibiotics | -662
supervening sepsis | -648
surgical treatment | -648
infected mesh removed | -648
open abdomen | -648
thick granulation tissue | -648
site of perforation confirmed | -648
Kehr drain | -648
vacuum-assisted system | -648
Negative Pressure Wound Treatment | -648
NPWT | -648
baby bottle nipple | -648
absorbable stitches | -648
biologic glue | -648
NPWT with low pressure | -648
stitches and glue dissolved | -636
unsuccessful efforts | -636
Hyalomatrix | -636
platelet gel | -636
non-cross-linked biologic implant | -636
biologic glue | -636
handmade “fistula patch” | -636
silastic drain | -636
fistula narrowed | -636
ECF | -636
catabolic status reversed | -636
antibiotics | -636
TPN | -636
improved general and local conditions | -120
surgery planned | -120
laparoscopic approach | -120
informed consent | -120
adhesiolysis | -120
laparotomy | -120
intestinal tract resection | -120
side to side jejuno-jejunostomy | -120
abdomen irrigated | -120
abdominal wall reconstructed | -120
anterior component separation | -120
absorbable mesh | -120
Prevena Incisional System | -120
postoperative course uneventful | -96
discharged | 16
follow-up | 1752
no complications | 1752
no hernia recurrence | 1752