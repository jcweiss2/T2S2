56 years old | 0
female | 0
anemia | 0
high sedimentation rate | 0
diabetes mellitus | -672
hypertension | -672
hyperthyroidism | -672
admitted to the hospital | 0
body temperature 38.0°C | 0
pulse rate 75 beats/min | 0
blood pressure 91/55 mm Hg | 0
tenderness on the left iliac fossa | 0
pleural effusions | 0
minimal infiltration | 0
levofloxacin IV 0.5 g antibiotic treatment | 0
blood and urine samples taken for culture | 0
Escherichia coli | 24
piperacillin/tazobactam and linezolid | 24
constipation | 72
diffuse distension and tenderness | 72
sluggish bowel sounds | 72
air-fluid levels | 72
free peritoneal fluid | 72
contrast-enhanced chest multidetector computed tomography (MDCT) scan | 72
bilateral pleural effusion | 72
compression atelectasis | 72
hypodense mass and calcifications at the right breast | 72
enlarged thyroid gland | 72
filling defect secondary to a free-floating thrombus | 72
partial obstruction of the descending thoracic aorta lumen | 72
massive ascites | 72
wedge-shaped renal infarction | 72
mild mitral regurgitation | 72
intravenous fluids | 72
broad spectrum antibiotics | 72
enoxaparin sodium | 72
total parenteral nutrition | 72
respiratory distress | 144
sepsis | 144
visceral ischemia | 144
transferred to the intensive care unit (ICU) | 144
unconscious | 168
intubated | 168
leukocyte count of 12.3×10^9 L | 168
hemoglobin levels of 10.5 g/dL | 168
thrombophilia workup was normal | 168
potassium 3.31 mmol/L | 168
creatinine 2.14 mg/dL | 168
lactate dehydrogenase 439 U/L | 168
albumin 2.79 g/dL | 168
emergency hemodialysis | 168
albumin replacement | 168
decrease in blood pressure | 168
positive inotropic agents | 168
cardiac arrest | 216
death | 216