33 years old | 0
    male | 0
    presented to the emergency department | 0
    fever | -24
    altered mental status | -24
    nausea | -48
    vomiting | -48
    diarrhea | -48
    visited emergency room | -48
    discharged to home | -48
    developed fever | 0
    became acutely confused | 0
    nonsensical speech | 0
    tonic clinic seizure | -24
    temperature of 39.1 °C | -24
    past medical history of HIV | -52704
    CD4+ cell count 1,782 cells/mm³ | -672
    HIV-1 RNA level < 20 copies/mL | -672
    antiretroviral therapy with DTG/3TC/ABC | -26208
    up-to-date vaccinations | -26208
    history of secondary syphilis | -26208
    presented with nasopharyngitis symptoms | -240
    Group A Streptococcus test negative | -240
    prescribed supportive care | -240
    temperature 39.1 °C | 0
    heart rate 114 beats/min | 0
    respiratory rate 32 breaths/min | 0
    blood pressure 163/94 mm Hg | 0
    oxygen saturation 100% | 0
    Glasgow Coma Scale score of 11 | 0
    nuchal rigidity | 0
    agitation | 0
    pupils equal and reactive | 0
    dental caries | 0
    clear pulmonary exam | 0
    lactic acid 14.79 mmol/L | 0
    sodium 143 mmol/L | 0
    potassium 3.1 mmol/L | 0
    chloride 109 mmol/L | 0
    CO2 12 mmol/L | 0
    BUN 14 mg/dL | 0
    creatinine 1.1 mg/dL | 0
    glucose 74 mg/dL | 0
    calcium 7.9 | 0
    anion gap 26 mmol/L | 0
    WBC 3.5 × 10³/µL | 0
    hemoglobin 12.7 g/dL | 0
    platelet 95 × 10³/µL | 0
    INR 1.6 | 0
    PT 18.9 s | 0
    alkaline phosphatase 226 IU/L | 0
    toxicology screen positive for marijuana | 0
    ethanol level < 10 mg/dL | 0
    CD4+ cell count 182 cells/mm³ | 0
    CT head unremarkable | 0
    blood cultures obtained | 0
    lumbar puncture performed | 0
    CSF yellow/turbid | 0
    CSF glucose < 10 mg/dL | 0
    CSF protein 1,185 mg/dL | 0
    CSF WBC 2,663/µL | 0
    cryptococcal antigen negative | 0
    VDRL test nonreactive | 0
    Gram smear of CSF with gram-negative diplococci | 0
    transferred to ICU | 0
    empiric vancomycin initiated | 0
    empiric ceftriaxone initiated | 0
    empiric ampicillin initiated | 0
    empiric acyclovir initiated | 0
    empiric dexamethasone initiated | 0
    intubated | 0
    sudden drop in blood pressure | 24
    PEA arrest | 24
    return of spontaneous circulation | 24
    required vasopressors | 24
    pupils dilated and non-reactive | 24
    CT head showed increased edema | 24
    unresponsive on physical exam | 24
    EEG suppression of activity | 24
    expired | 48
    blood cultures positive for H. influenzae | 48
    CSF cultures positive for H. influenzae | 48
    NTHi biotype I | 48
    cause of death sepsis | 48
    cause of death meningitis | 48
<|eot_id|>
