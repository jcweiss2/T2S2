66 years old | 0 | 0 
male | 0 | 0 
dual-chamber pacemaker | -10512 | -10512 
sick sinus syndrome | -10512 | -10512 
paroxysmal atrial fibrillation | -10512 | -10512 
severe lumbar back pain | -24 | 0 
mental status changes | -12 | 0 
hypotension | -12 | 0 
acute renal failure | -12 | 0 
hypoxemic respiratory failure | -12 | 0 
emergent intubation | -12 | 0 
severe sepsis | -12 | 0 
hemodynamic support | -12 | 0 
vasopressin | -12 | 0 
norepinephrine | -12 | 0 
blood cultures | -12 | 0 
methicillin-sensitive Staphylococcus aureus | -12 | 0 
vancomycin | -12 | -6 
nafcillin | -6 | 0 
transthoracic echocardiogram | -6 | 0 
left ventricular ejection fraction | -6 | 0 
patent foramen ovale | -6 | 0 
computed tomography scan | -6 | 0 
osteomyelitis | -6 | 0 
magnetic resonance imaging | -6 | 0 
septic emboli | -6 | 0 
transesophageal echocardiogram | -6 | 0 
vegetation | -6 | 0 
pacemaker lead | -6 | 0 
tricuspid valve | -6 | 0 
right ventricle | -6 | 0 
cardiothoracic surgery | -6 | 0 
laser lead extraction | 0 | 72 
Indigo Penumbra system | 0 | 72 
intracardiac echocardiography | 0 | 72 
aspiration | 0 | 72 
vegetation removal | 0 | 72 
RA lead extraction | 72 | 72 
RV lead extraction | 72 | 72 
pathology | 72 | 72 
gram-positive cocci | 72 | 72 
methicillin-sensitive Staphylococcus aureus | 72 | 72 
condition improved | 0 | 48 
condition worsened | 72 | 96 
tissue necrosis | 96 | 96 
lactic acidosis | 96 | 96 
renal failure | 96 | 96 
care withdrawn | 96 | 96 
extubation | 96 | 96 
death | 96 | 96