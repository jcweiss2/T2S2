44 years old | 0
man | 0
rash on left forehead | -72
vesicle on left forehead | -72
headache | -144
fever (38°C and higher) | -72
diagnosed with HZO | -72
antiviral drugs | -72
analgesics | -72
hospitalized | -72
worsening left-sided frontal headache | 0
nausea | 0
blurred vision | 0
diplopia | 0
transferred to hospital | 0
alert | 0
febrile (38.3°C) | 0
crust on forehead | 0
normal cardiopulmonary findings | 0
normal neurological findings | 0
heart rate 78 beats/min | 0
blood pressure 110/60 mmHg | 0
respiratory rate 20 breaths/min | 0
visual acuity 6/12 bilaterally | 0
no ocular tissue abnormalities | 0
no visual field defects | 0
horizontal diplopia | 0
lateral rectus muscle paresis | 0
6th cranial nerve palsy | 0
no facial infection | 0
no periorbital swelling | 0
no respiratory tract infection | 0
no urinary tract infection | 0
no skin infection | 0
WBC count 10,100 mm3 | 0
elevated erythrocyte sedimentation rate (120 mm/h) | 0
elevated C-reactive protein (10.17 mg/dl) | 0
blood culture | 0
no CSF analysis | 0
MRI showing cavernous sinus thrombosis | 0
superior ophthalmic vein thrombosis | 0
admitted to ICU | 0
neurologist consultation | 0
infectious medicine consultation | 0
no diabetes mellitus | 0
no hypertension | 0
dental treatment 3 months ago | -2160
left maxillary pain 1 month ago | -720
antibiotic treatment | 0
second-generation cephalosporin | 0
Streptococcus constellatus in blood culture | 0
switched to clindamycin | 0
echocardiography performed | 0
no infective endocarditis | 0
low molecular weight heparin | 0
improved symptoms after 7 days | 168
discharged | 168
no complications during follow-up | 168
