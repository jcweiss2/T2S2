50 years old | 0
male | 0
admitted to the hospital | 0
progressive dyspnea | -168
cough | -168
cold sweats | -168
night sweating | -8760
weight loss | -8760
HIV infection | -104544
double-sided pneumonia | -168
Pneumocystis jirovecii | -168
acquired immunodeficiency syndrome (AIDS) | -168
antiretroviral therapy | -104544
undetectable viral load | -8760
stopped taking medication | -8760
lived in a homeless shelter | -8760
no intravenous drug use | 0
no alcohol use | 0
quit smoking | -131040
physical examination | 0
tachypneic | 0
oxygen saturation 88% | 0
blood pressure 130/80 mmHg | 0
heart rate 132 per minute | 0
temperature 38.2°C | 0
percussion of the lungs | 0
auscultation | 0
normal breath sounds | 0
hemoglobin 7.2 mmol/L | 0
white blood cell count 6.6 × 10^9/L | 0
platelets 214 × 10^9/L | 0
C-reactive protein (CRP) 64 mg/L | 0
no renal or hepatic insufficiency | 0
CD4: 0.039 × 10^9/L | 0
CD8: 1.2 × 10^9/L | 0
CD4/CD8 ratio: 0.033 | 0
chest X-ray | 0
bilateral cloudy infiltrates | 0
treated according to the local sepsis protocol | 0
gentamicin 280 mg | 0
amoxicillin/clavulanic acid 1200 mg | 0
cotrimoxazole (3 × 1920 mg) | 24
prednisolone (2 × 40 mg) | 24
bronchoscopy with bronchoalveolar lavage (BAL) | 48
dyspneic | 48
low oxygen saturations (82%) | 48
subcutaneous emphysema | 48
endotracheal intubation | 48
mechanical ventilation | 48
computed tomography (CT) scan of the chest | 48
subcutaneous and mediastinal emphysema | 48
severe air bronchograms | 48
bilateral infiltrations | 48
admitted to the intensive care unit (ICU) | 48
increased subcutaneous and mediastinal emphysema | 72
swelling of the entire face, arms, and torso | 72
several bronchoscopies | 72
no tracheal injury | 72
lung protective ventilation | 72
low tidal volumes | 72
low airway pressures | 72
new CT scan | 168
severe subcutaneous and mediastinal emphysema | 168
treatment of the emphysema by skin incisions | 168
fear of viral spreading | 168
VAC therapy | 216
infraclavicular skin incisions | 216
improvement of subcutaneous emphysema | 216
gradual clinical improvement | 216
VAC therapy ended | 225
subcutaneous emphysema continued to decrease | 225
inflammatory markers decreased | 216
pulmonary infiltrations on the chest X-ray decreased | 216
adequate treatment of the PJP | 216
extubated | 408
ICU-acquired weakness | 408
dysphonia | 408
discharged to the general ward | 600
antiretroviral medicine restarted | 600
discharged to a medical rehabilitation center | 720