26 6/7 weeks gestational age | 0
female | 0
admitted to the Neonatal Intensive Care Unit | 0
prematurity | 0
respiratory distress syndrome | 0
chronic lung disease | 0
suspected sepsis | 0
metabolic acidosis | 0
anemia | 0
suspected necrotizing enterocolitis | 0
cow’s milk protein allergy | 0
diagnosis of SCD | 10
SCD-SS type | 5
irritable | 83
swelling of the left thigh | 83
tenderness | 83
minimal active movement | 83
non-displaced fracture of the left femoral shaft | 83
periosteal reaction | 83
splint placed | 83
healing fracture | 93
calcium normal | 83
phosphorus normal | 83
vitamin D normal | 83
alkaline phosphatase level 599 units/L | 79
alkaline phosphatase level peak 699 units/L | 14
vitamin D supplementation added | 83
bluish sclera | 83
diagnosis of OI type 1 | 83
13th percentile for length | 18
below third percentile for weight | 18
no further fractures | 18
hospitalized for sickle cell pain crises (age 1 year) | 12
irritable (age 1 year) | 12
inability to bear weight on right lower extremity (age 1 year) | 12
imaging no new fractures (age 1 year) | 12
hospitalized for sickle cell pain crises (age 16 months) | 16
irritable (age 16 months) | 16
inability to bear weight on right lower extremity (age 16 months) | 16
imaging no new fractures (age 16 months) | 16
folic acid | 18
prophylactic penicillin | 18
vitamin D supplementation | 18
blue sclera | 18
height 13th percentile | 18
weight below third percentile | 18
referred to comprehensive center for OI | 18
