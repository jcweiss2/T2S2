39 years old|0
    male|0
    admitted to the emergency department|0
    paraesthesia in all limbs| -48
    diplopia| -48
    nausea| -48
    weakness in both lower limbs|0
    weakness in both upper limbs|0
    bilateral abducens nerve paralysis|0
    facial diplegia|0
    flaccid areflexic paralysis of the limbs|0
    Medical Research Council grade 3/5 in all muscles of the upper extremities|0
    Medical Research Council grade 2/5 in lower extremities|0
    bilateral flexor plantar responses|0
    bowel not involved|0
    bladder not involved|0
    electromyography examination|0
    acute, acquired, disseminated polyneuropathy syndrome|0
    prolongation of the distal motor latency|0
    prolongation of the F-wave|0
    decreased sensory nerve amplitude|0
    decreased motor nerve amplitude|0
    disperse responses|0
    reduced nerve conduction velocities|0
    cerebrospinal fluid elevated protein concentration|0
    cerebrospinal fluid normal cell count|0
    anti-ganglioside antibodies negative|0
    intravenous immune globulin (IVIG) administrated|0
    weakness progressed rapidly|24
    unable to stand|24
    6th cranial nerve involvement|24
    7th cranial nerve involvement|24
    respiratory muscle weakness|24
    respiratory failure|24
    mechanical ventilation|24
    remained in the intensive care unit for two months|0
    IVIG administrated again over 5 days| -48
    plasmapheresis performed on every other day| -48
    booster IVIG continued every 15 days| -48
    rehabilitation performed from the beginning of the disease|0
    oral prednisolone administered|0
    prednisolone reduced by 5 mg every two weeks|0
    pain in both hips| -1344
    decreased range of motion (ROM) in both hips| -1344
    NHO diagnosed| -1344
    serum calcium 10.5 mEq/L| -1344
    serum alkaline phosphatase 61 IU/L| -1344
    intravenous ibandronic acid given weekly| -1344
    IV ibandronic acid discontinued| -1344
    etidronate disodium administered| -1344
    ALP levels measured periodically| -1344
    Ca levels measured periodically| -1344
    rehabilitative management continued| -1344
    passive ROM exercises| -1344
    active - assistive ROM exercises| -1344
    breathing exercises| -1344
    electrotherapy| -1344
    discharged from the ICU| -1344
    muscle strengths improved in upper extremities| -1344
    muscle strengths improved in lower extremities| -1344
    stand up with support| -1344
    cannot walk| -1344
    cannot sit in low position| -1344
    passive ROM of both hips restricted| -1344
    three-phase bone scan study showed Tc99m-MDP uptake| -1344
    computed tomography guidance| -1344
    corticosteroid injection made| -1344
    pain decreased| -1344
    10º degree flexion achieved| -1344
    rehabilitation program continues| -1344
    walk with a walker| -1344
    sit without support| -1344
    <|eot_id|>
    