49 years old | 0
male | 0
admitted to emergency department | 0
worsening fever | -168
cough | -168
shortness of breath | -168
febrile | 0
tachycardic | 0
hypoxic | 0
SpO2 of 70% | 0
nasal cannula oxygen supplementation | 0
SpO2 improved to 92%-95% | 0
white blood cell count of 11.3 × 10^9/L | 0
lactate dehydrogenase of 3,147 units/L | 0
C-reactive protein of 265.9 mg/L | 0
ferritin of 1,760 ng/mL | 0
D-dimer of 124,802 ng/mL | 0
acute hypoxic respiratory failure | 0
COVID-19 virus infection | 0
real-time reverse transcriptase polymerase chain reaction test for SARS-CoV-2 RNA | 0
positive SARS-CoV-2 RNA | 0
empiric antibiotics with ceftriaxone and azithromycin | 0
low-weight-molecular heparin therapy with enoxaparin | 0
steroid course with dexamethasone | 0
antiviral therapy with remdesivir | 0
convalescent plasma therapy refused | 0
inflammatory markers increased | 24
tocilizumab | 24
dyspneic | 336
exercise in room | 336
nonrebreather mask | 336
oxygen 10-15 L/min | 336
large right pneumothorax | 336
mediastinal shift | 336
CT-guided chest tube placement | 336
8.5-French pigtail catheter | 336
low intermittent suction | 336
persistent right pneumothorax | 336
second 22-French chest tube | 336
mildly improved right pneumothorax | 336
transferred to intensive care unit | 336
worsening respiratory status | 336
antibiotic therapy broadened | 336
immunosuppressive therapy continued | 336
dexamethasone | 336
chest tube advanced to 36-French size | 336
large air-filled bullous process | 336
suspicious for bronchopulmonary fistula | 336
intubated | 336
impending respiratory failure | 336
cardiothoracic surgery consulted | 336
right middle invasive thoracotomy | 336
right bronchopleural fistula repair | 336
pleurodesis | 336
large bronchopleural fistula | 336
necrotic empyema | 336
repaired | 336
resected | 336
intraoperative specimens sent for pathological evaluation | 336
initial cultures concerning for fungal process | 336
probable mucormycosis | 336
amphotericin B | 336
worsening respiratory failure | 504
septic shock | 504
maximum vasopressor and antimicrobial therapy | 504
marked bradycardia | 504
asystole | 504
expired | 504
microbiological analysis of intraoperative specimens | 508
positive for Rhizopus species | 508