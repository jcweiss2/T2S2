55 years old | 0
male | 0
multiple myeloma | -672
previous stem cell transplant | -672
recurrence of disease | -672
carfilzomib treatment | -48
fever | -48
dyspnea | -72
productive cough | -72
admitted to the hospital | 0
febrile | 0
tachypneic | 0
tachycardic | 0
alert and fully oriented | 0
normal blood pressure | 0
decreased breath sounds in the right lung base | 0
pancytopenia | 0
white blood cell count of 1.2 × 109/l | 0
hemoglobin of 53 g/l | 0
platelets of 4.0 × 109/l | 0
treated with cefepime and azithromycin | 0
acyclovir treatment | 0
allopurinol treatment | 0
fluconazole treatment | 0
pantoprazole treatment | 0
new-onset hypoxia | 2
hypotension | 2
altered mental status | 2
transferred to the medical intensive care unit | 2
lactic acid of 6.1 mMol/l | 2
pH of 7.40 | 2
carbon dioxide partial pressure (PaCO2) of 3.3 kPa | 2
PaO2 of 11.3 kPa | 2
measured O2sat of 94% | 2
intubation procedure | 2
treated with topical endobronchial lidocaine | 2
intravenous etomidate | 2
succinylcholine | 2
increasingly hypoxic | 4
brownish arterial blood gas (ABG) | 4
pH of 7.21 | 4
PaCO2 of 3.3 kPa | 4
PaO2 of 55.1 kPa | 4
measured O2sat of 49% | 4
co-oximetry | 4
methemoglobin level of 53% | 4
intravenous methylthioninium chloride | 4
methemoglobin level of 12% | 4.5
methemoglobin level of 9% | 5
O2sat > 90% | 5
bright red coloration to the ABG sample | 5
septic shock | 24
bacteremia with Rothia mucilaginosa | 24
death | 48