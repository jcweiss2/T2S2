19 years old | 0
male | 0
admitted to the hospital | 0
meningococcal meningitis | 0
multi-organ failure | 0
acute renal insufficiency | 0
amputation of the right lower leg | 0
neurological sequelae | 0
prolonged immobilization | 0
hypercalcaemia | -1440
maximum corrected serum calcium concentration of 3.4 mmol/L | -1440
serum parathyroid hormone (PTH) concentration was below the detection limit | -1440
immobilization-related hypercalcaemia | -1440
pamidronate | -720
near normalization of the serum calcium concentration | -720
increased serum calcium concentration | -480
pamidronate | -480
near-normal level of serum calcium concentration | -480
renal function remained stable | -480
high serum phosphate level | -480
discharged to a rehabilitation centre | -480
mobilization was limited | -480
persistent renal insufficiency | -480
eGFR of 24 mL/min/1.73 m² | -480
increased serum calcium concentration | 0
nausea | 0
vomiting | 0
readmitted to the hospital | 0
hyperhydration | 0
oral furosemide | 0
calcitonin | 0
decreased serum calcium concentration | 24
low serum 25-OH-vitamin D | 24
low serum 1,25-di-OH-vitamin D | 24
no PTH-related peptide | 24
high urinary calcium excretion | 24
normal urinary metanephrines | 24
normal serum thyroid stimulating hormone | 24
normal cortisol | 24
normal aluminium concentrations | 24
normal free light chain kappa/lambda ratio | 24
no lymphadenopathy | 24
no skeletal metastasis | 24
denosumab | 168
decreased serum calcium concentration | 168
decreased serum phosphate level | 168
effective inhibition of bone resorption | 168
supplementation with calcium-carbonate/colecalciferol and active vitamin D | 168
normalized serum calcium concentration | 168
increased serum PTH concentration | 168
normal serum calcium concentration | 336
stopped vitamin D and calcium supplementation | 336