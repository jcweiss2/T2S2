27 years old | 0
woman | 0
transferred to our department | 0
seizure episodes | -24
loss of consciousness | -24
admitted to a local psychiatric department | -72
acute psychosis | -72
spoke few words | -72
restless | -72
unwilling to eat | -72
cold-like symptoms | -168
runny nose | -168
low-grade fever | -168
physical examination | 0
vital signs stable | 0
body weight 52.0 kg | 0
height 163 cm | 0
neurological examination | 0
Glasgow coma scale score 6 | 0
Eye opening 1 | 0
Verbal response 1 | 0
Motor response 4 | 0
laboratory results not remarkable | 0
electroencephalogram results not remarkable | 0
cranial magnetic resonance imaging | 0
mild signal changes bilateral hippocampus | 0
mild signal changes left temporal cortex | 0
local meningeal congestion | 0
anti-NMDA receptor antibodies detected | 0
serum anti-NMDA receptor antibodies 1:1000 | 0
cerebrospinal fluid anti-NMDA receptor antibodies 1:100 | 0
abdominal ultrasound screening | 0
weak liquid echo right ovary | 0
teratoma suspected | 0
tumor removal initiated | 24
pathology confirmed teratoma | 24
comatose | 0
persistent facial involuntary movement | 0
lip perastalsis | 0
uncontrolled eye blinking | 0
treated with large dose anesthetic agents | 0
diagnosis of anti-NMDA receptor encephalitis | 0
first-line therapy | 24
intravenous methylprednisolone pulse | 24
intravenous immunoglobin | 24
plasmapheresis | 24
immunoadsorption | 24
refractory to treatments | 24
neurological status not improve | 24
high anti-NMDA receptor antibody titers | 24
second-line therapy | 168
rituximab | 168
intravenous cyclophosphamide | 168
no reaction to second-line therapy | 168
bilateral salpingo-oophorectomy | 1272
inflammation observed | 1272
no teratoma observed | 1272
immunosuppressant therapy | 1272
mycophenolate mofetil | 1272
intrathecal methotrexate | 1272
intrathecal dexamethasone | 1272
antibody titer in CSF decreased | 1272
antibody titer 1:10 | 1464
awoke after 17 months | 1464
Glasgow coma scale score 9T | 1464
open and close eyes | 1464
extend tongue | 1464
turn head | 1464
physical therapy | 2928
good prognosis | 2928
mRS score 1 | 2928
diffuse muscular ossification | 2928
septicemia with Staphylococcus caprae | 552
septicemia with Klebsiella pneumoniae | 1968
heterotopic ossification | 2928
