32 years old | 0
female | 0
Indigenous | 0
G5T2A2L2 | 0
admitted to the hospital | 0
opioid withdrawal | -72
anemia | -72
malnourishment | -72
hypertension | -72
severe edema | -72
sepsis | -72
5 years of opioid intravenous drug use | -7200
2 g/d of fentanyl | -7200
0.5 g/d methamphetamine | -7200
10 cigarettes daily | -7200
previous hospital admissions | -7200
methadone | -7200
slow-release oral morphine | -7200
oral hydromorphone | -7200
iOAT offered | -7200
sepsis | -7200
IVDU | -7200
endocarditis | -7200
sublingual buprenorphine | -7200
precipitated withdrawal | -7200
adverse reactions | -7200
buprenorphine subcutaneous extended release | -7200
teratogenicity | -7200
community prenatal care | -7200
stable housing | 0
income assistance | 0
partner | 0
biological father | 0
IV fentanyl | -1
caesarean section | 0
APGARS of 6, 8, and 9 | 0
postpartum hemorrhage | 0
intrauterine balloon tamponade | 0
blood transfusion | 0
anesthesia support | 0
iOAT | 0
Pasero Opioid-induced Sedation Scale | 0
20 mg IV hydromorphone | 0
120 mg three times a day | 24
32 mg every hour | 24
70 mg oral methadone | 24
highest dose of iOAT | 120
120 mg IV hydromorphone | 120
60 mg q1h PRN oral hydromorphone | 120
100 mg oral methadone | 120
infant admitted to NICU | 0
respiratory distress | 0
meconium aspirations | 0
NICU | 0
ESC model | 0
nasogastric feeds | 24
0.04 mg/kg q4h PRN oral morphine | 48
0.12 mg q4h and 0.06 mg q4h PRN oral morphine | 144
maximum weight loss 5.8% | 144
infant transferred from NICU to FIR | 144
informed consent discussion | 0
breastfeeding on iOAT | 216
maternal HIV PCR test | 216
96 hours substance-free | 216
transfer to mother-infant rooming-in unit | 216
48-hour minimum observation period | 216
infant’s morphine discontinued | 216
morphine PRN ordered | 216
72 mL expressed breast milk | 216
110 mg IV hydromorphone BID | 216
155 mL of formula | 240
0.10 mg q4h PRN of morphine | 240
110 mg IV hydromorphone | 240
infant latched to breast | 240
infant monitored for NAS symptoms | 240
no clinically relevant apneas | 240
no bradycardias | 240
no desaturations | 240
no signs of respiratory depression | 240
no excessive sedation | 240
cardiopulmonary monitoring | 240
oxygen saturation | 240
q1h vitals | 240
q3h vitals | 240
337 mL EBM | 264
385 mL of formula | 264
no breastfeeding | 264
one low respiratory rate of 28 bpm | 264
saturation was 100% | 264
ESC reassuring | 264
340 mL EBM | 288
440 mL formula | 288
infant latched to breast for 30 minutes | 288
off morphine | 288
gaining weight | 288
no symptoms of sedation | 288
no respiratory depression | 288
no NAS | 288
transferred back to FIR | 288
mixed feeds | 288
maternal iOAT titrated down | 288
methadone titrated up | 288
addition of slow-release oral morphine | 288
discharged | 1104
190 mg methadone | 1104
1200 mg slow-release oral morphine | 1104
no evidence of maternal substance use | 1104
voluntary urine drug screens | 1104
Ages & Stages Questionnaire | 1248
infant scored above the cutoff score | 1248
communication | 1248
gross motor | 1248
fine motor | 1248
problem solving | 1248
personal-social | 1248
regained custody of her two other children | 1248