50 years old| 0
    man | 0
    alcoholism | 0
    admitted to an emergency hospital | 0
    worsening pain | -48
    redness of the right elbow | -48
    trivial trauma | -48
    X-ray of the elbow negative | 0
    discharged | 0
    non-steroidal anti-inflammatory drugs (NSAIDs) | 0
    persistent erythema | 24
    tenderness around his elbow | 24
    no systemic inflammatory symptoms | 24
    skin erythema | 24
    edema | 24
    warmness | 24
    tenderness on the right elbow | 24
    no axillar lymphadenopathy | 24
    white blood cell count of 7770/μL | 24
    CRP 533.6 mg/L | 24
    hemoglobin 14.8 g/dL | 24
    glucose 0.83 g/L | 24
    creatine 1.4 mg/dL | 24
    sodium 133 mmol/L | 24
    LRINEC score of 6 | 24
    kidney function tests normal | 24
    liver function tests normal | 24
    blood culture negative | 24
    diagnose of cellulitis | 24
    intravenous antibiotics (Cefazoline 4 g daily and Metronidazole 1500 mg daily) | 24
    condition continued to deteriorate | 168
    intense pain | 168
    significant edema | 168
    tenderness of his right elbow | 168
    wound culture revealed Streptococcus pyogenes infection | 168
    brought to our hospital | 168
    febrile (38°C) | 168
    blood pressure 148/83 mmHg | 168
    white blood cell count of 16000/μL | 168
    CRP 95 mg/L | 168
    LRINEC score of 3 | 168
    blood endotoxin negative | 168
    margins of tenderness spread all over the right upper extremity | 168
    erythema spread all over the right upper extremity | 168
    upper right thorax with phlyctens | 168
    areas of necrosis | 168
    emergency aggressive debridement of necrotic tissues | 168
    general anesthesia | 168
    skin swabs taken during the operation negative | 168
    underlying muscles intact | 168
    transferred to the intensive care unit | 168
    respiratory support | 168
    renal support | 168
    circulatory support | 168
    intensive debridement | 168
    intravenous penicillin (4.000.000 UI, 6 times daily) | 168
    multiple sets of vacuum-assisted closure (VAC) technique | 168
    hyperbaric oxygen therapy (HBOT) | 168
    wound closed by split-thick-ness skin graft | 408
    no complications | 408
    discharged | 432
    totally healed wounds | 432
    stiff elbow | 432
    regained an acceptable range of motion of his right arm | 1752
    no sign of infection recurrence | 17520
    