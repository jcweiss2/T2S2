53 years old | 0
    female | 0
    myeloablative allogeneic hematopoietic cell transplant | -9504
    relapsing acute lymphoblastic leukaemia | -9504
    relapse after BMT | -9504
    CAR-T therapy targeting CD19 | -9504
    cyclophosphamide | -9504
    fludarabine | -9504
    grade 1 cytokine release syndrome (CRS) | -9504
    tocilizumab | -9504
    methylprednisolone 50 mg | -9504
    prophylactic levetiracetam | -9504
    stopped levetiracetam | -9504
    improved neurotoxicity (confusion) | -9504
    admitted to the ward | 0
    ongoing pancytopenia | 0
    fevers | 0
    Escherichia coli bacteraemia | 0
    treated bacteraemia | 0
    new fevers | 0
    dyspnoea | 0
    hypoxemia | 0
    requiring 2 L continuous oxygen | 0
    chest CT consolidations | 0
    vancomycin-resistant enterococcal bacteraemia | 0
    prophylactic foscarnet | 0
    prophylactic pentamidine | 0
    prophylactic isavuconazole | 0
    prophylactic levofloxacin | 0
    broadened meropenem | 0
    broadened linezolid | 0
    restlessness | 0
    agitation | 0
    obtundation | 0
    intubation | 0
    ICU transfer | 0
    normal basic metabolic panel | 0
    mild elevation of total bilirubin | 0
    minor increased INR | 0
    malnutrition | 0
    normal kidney function | 0
    normal BUN level | 0
    ongoing pancytopenia | 0
    WBC 0.0×10^9/L | 0
    hemoglobin 6.7 g/dL | 0
    platelet count 16×10^9/L | 0
    encephalopathy workup | 0
    normal thyroid-stimulating hormone | 0
    normal vitamin B1 | 0
    normal vitamin B12 | 0
    negative electroencephalogram | 0
    negative head CT | 0
    lumbar puncture | 0
    0 WBC in CSF | 0
    0 RBC in CSF | 0
    protein 21 mg/dL | 0
    glucose level 82 mg/dL | 0
    negative gram stain | 0
    negative bacterial culture | 0
    negative fungal culture | 0
    negative herpes simplex virus PCR | 0
    negative cytomegalovirus PCR | 0
    negative varicella zoster virus PCR | 0
    negative cryptococcal antigen | 0
    negative cytology | 0
    negative flow analysis | 0
    ammonia level 391 µmol/L | 0
    CT abdomen and pelvis | 0
    ultrasound abdomen | 0
    anasarca | 0
    hypoalbuminaemia | 0
    doxycycline added | 0
    oral lactulose | 0
    methylprednisolone 1 g/day | 0
    bronchoscopy with BAL | 0
    BAL bacterial culture | 0
    BAL fungal culture | 0
    BAL viral PCR | 0
    BAL Ureaplasma PCR | 0
    ammonia level 643 µmol/L | 24
    epileptiform activity | 24
    high-dose benzodiazepine infusion | 24
    levetiracetam | 24
    lacosamide | 24
    propofol infusion | 24
    pentobarbital initiated | 24
    halted status epilepticus | 24
    CT head mild cerebral oedema | 24
    renal replacement therapy | 24
    ammonia level 258 µmol/L | 24
    changed meropenem to ceftazidime/avibactam | 24
    added amphotericin B | 24
    added acyclovir | 24
    genetics consult | 48
    hyperammonemia assessment | 48
    negative urine organic acids | 48
    negative urine orotic acid | 48
    negative plasma amino acids | 48
    negative plasma acylcarnitine | 48
    negative genetics testing | 48
    dextrose 10% infusion | 48
    levocarnitine | 48
    arginine infusion | 48
    sodium phenylbutyrate | 48
    ammonia levels 270 µmol/L | 48
    MRI brain diffuse cerebral oedema | 72
    positive Ureaplasma PCR | 72
    added levofloxacin | 72
    progression in brain damage | 72
    family elected to withdraw care | 72
    patient died | 72
    
    
    <|end_header_id|>

