Here is the table of events and timestamps:

age | 0
sex | 0
male | 0
65 years old | 0
presented to the emergency | 0
multiple blisters and erosions | 0
oral mucosa | 0
scalp | 0
maggot infection | 0
previous episodes of lesions | -6 months
previous treatment with steroids and generic medications | -12 months
developed lesions | -6 months
worsened | -6 months
febrile | 0
Nikolsky sign | 0
positive | 0
diagnosis of PV | 0
skin biopsy | 0
tzanck smear | 0
intravenous dexamethasone pulse | 0
fluids | 0
fresh frozen plasma | 0
dressings | 0
intravenous antibiotics | 0
Piperacillin/Tazobactam | 0
Teicoplanin | 0
pus culture and sensitivity | 0
adjuvant immunosuppressors | 0
held back | 0
infection | 0
shifted to ICU | 0
oozing from skin ulcerations | 0
hemorrage excoriation with peeling of skin | 0
oral methyl prednisolone | 0
no improvement | 0
general condition worsened | 0
hypoproteinemia | 0
pleural effusion | 7
enterobacter | 7
Staphylococcus aureus | 7
Proteus mirabilis | 7
intravenous Tigecycline | 7
vancomycin | 7
erosions persisted | 7
new blisters | 7
sepsis | 7
high grade fever | 7
albumin levels fell | 7
TPE cycle | 7
plasma exchange | 7
intermittent cell separator | 7
femoral access | 7
12-French double lumen dialysis catheter | 7
citrate | 7
isotonic sterile saline | 7
4% purified human albumin | 7
FFP | 7
hemodynamic parameters | 7
complications | 7
calcium gluconate | 7
hemogram | 7
serum electrolytes | 7
total protein | 7
albumin | 7
Nikolsky sign became negative | 7
no new lesions | 7
exudation from lesions reduced | 7
dressings remained dry | 7
re-epithelization | 7
healing | 7
oral lesions healed | 7
little erosions persisted | 7
pulse therapy of IV methyl prednisolone | 7
cyclophosphamide | 7
further improvement | 7
clinically stable | 7
another TPE cycle | 7
cost restraint | 7
discharged | 7
maintained dose of IV dexamethosone pulse | 7
daily oral prednisolone | 7