72 years old | 0
male | 0
pulmonary fibrosis | 0
oral steroids | 0
home oxygen therapy | 0
hypertension | 0
diabetes mellitus | 0
no prior smoking history | 0
progressive dyspnea | -504
cough | -504
yellow sputum | -504
no hemoptysis | -504
fever | -168
night sweats | -168
six-pound weight loss | -168
rapidly growing scalp lesion | -1344
pain | -1344
no pruritus | -1344
no discharge | -1344
denied exposure to smoke | 0
denied tuberculosis exposure | 0
temperature 96.8°F | 0
blood pressure 153/87 | 0
heart rate 82 | 0
respiratory rate 22 | 0
oxygen saturation 86% | 0
large ulcerative scalp lesion | 0
no cervical lymphadenopathy | 0
bilateral diffuse crackles | 0
leukocytosis | 0
white blood count 23,200 Cells/mcL | 0
hemoglobin 12.3 g/dL | 0
platelets 211,000/mcL | 0
blood urea nitrogen 17 mg/dL | 0
creatinine 0.8 mg/dL |. 0
arterial blood gas pH 7.44 | 0
PO2 51 | 0
PCO2 39 | 0
chest X-ray bilateral interstitial infiltrates | 0
admitted to medical floor | 0
intravenous corticosteroids | 0
oxygen | 0
nebulized treatments | 0
symptomatic improvement | 0
echocardiogram severe pulmonary hypertension | 0
CT chest diffuse fibrotic changes | 0
multiple densities | 0
CT-guided lung biopsy | 0
poorly differentiated malignant neoplasm | 0
necrosis | 0
immunohistochemical stains adenocarcinoma | 0
EGFR negative | 0
RAS negative | 0
alk translocation negative | 0
scalp lesion excision | 0
pathology poorly differentiated adenocarcinoma | 0
immunohistochemical confirmation | 0
severe hypoxic respiratory failure | 0
intubation | 0
transfer to ICU | 0
septic shock | 0
healthcare-associated pneumonia | 0
vasopressors | 0
intravenous antibiotics | 0
poor prognosis | 0
condition deteriorated | 0
expired | 336
