term male neonate | 0
born by normal spontaneous vaginal delivery | 0
mom with normal prenatal screens | -672
gestational diabetes | -672
hydronephrosis with stent placement | -672
multiple urinary tract infections secondary to Klebsiella sp | -672
membranes spontaneously ruptured for 13 h with clear fluid | -13
temperature instability | 0
respiratory distress with increasing supplemental oxygen requirement | 0
transferred to the neonatal intensive care unit (ICU) | 0
dusky with oxygen saturations of 80% | 0
placed on 2 L of nasal cannula at 21% FiO2 | 0
continued to exhibit signs of respiratory distress including grunting and tachypnea | 0
FiO2 was increased to 40% | 0
improved | 0
serum glucose, blood gas, complete blood count, renal function panel, and C-reactive protein were unremarkable | 0
chest radiograph showed mild diffuse ground glass opacities without focal consolidation | 0
blood culture was drawn | 0
empirically started on ampicillin, gentamicin, and ceftazidime | 0
respiratory failure on day 2 of admission | 48
intubation | 48
copious purulent drainage from his left eye | 48
ophthalmologic examination revealed diffuse fleshy red pseudomembrane coating the bulbar and tarsal conjunctiva of the left eye | 48
pseudomembrane coating was debrided yielding purulent and serosanginous drainage | 48
bacterial culture from the left eye grew pan-sensitive E. coli | 48
viral culture did not demonstrate any growth | 48
blood and urine cultures did not demonstrate any growth | 48
cerebral spinal fluid studies were collected | 48
cerebral spinal fluid studies were negative | 48
mom’s placental pathology did not show any abnormal findings | 0
patient’s mother was hospitalized shortly after delivery for urosepsis secondary to E. coli | 0
sensitivities of E. coli recovered from the mother’s urine culture mirrored that of the infant’s E. coli isolated from his ocular drainage | 0
successfully extubated to nasal cannula | 72
repeat ophthalmologic examinations showed significant clinical improvement after 24–48 h of intravenous and topical antimicrobials | 72
completed a full 14-day course of antimicrobial therapy with ampicillin | 168
completed 11 days of moxifloxacin eye drops | 168
weaned to room air on day of life 5 | 120
ready to be discharged home when the antibiotic course was complete | 168
follow-up eye examination 1 week after discharge was normal | 216
showing complete resolution of conjunctivitis | 216