3 years old | 0
male | 0
admitted to the hospital | 0
cough | -48
cold | -48
fever | -48
poor oral intake | -48
febrile convulsions | -720
vomiting | -720
cyanosis | -720
deviation of eyes | -720
loss of consciousness | -720
electroencephalogram | -720
cerebrospinal fluid studies | -720
neuroimaging | -720
atypical febrile convulsions | -720
birth history normal | 0
developmental history normal | 0
no family history of epilepsy | 0
febrile | 0
mild congestion in the throat | 0
symptomatic treatment | 0
high-grade fever | 4
vomiting | 4
bluish discoloration of the extremities | 4
tachypnea | 4
deviation of both eyes to the right side | 4
unresponsive | 4
loose stools | 4
drowsy | 4
temperature 39.9°C | 4
oxygen saturation 90% | 4
blood pressure 72/30 mmHg | 4
respiratory rate 39/min | 4
heart rate 220/min | 4
fluid resuscitation | 4
high flow oxygen | 4
phenytoin | 4
sinus tachycardia | 4
shifted to Intensive Care Unit | 4
regaining consciousness | 6
hemodynamically stable | 6
fully conscious | 9
normal neurological examination | 24
discharged | 72
phenytoin stopped | 96
asymptomatic | 1488
normal neurological examination | 1488
normal neuroimaging | 1488
normal EEG | 1488