83 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
admitted to the hospital | 0 | 0 | Factual
syncope | -24 | -24 | Factual
fell to the ground | -24 | -24 | Factual
leg ecchymosis | 0 | 0 | Factual
anuric | 0 | 0 | Factual
rhabdomyolysis-induced AKI | 0 | 0 | Factual
sepsis | 0 | 0 | Factual
acute prostatitis | 0 | 0 | Factual
increased urea | 0 | 0 | Factual
increased creatinine | 0 | 0 | Factual
increased myoglobin | 0 | 0 | Factual
increased CPK | 0 | 0 | Factual
increased LDH | 0 | 0 | Factual
increased CRP | 0 | 0 | Factual
increased PCT | 0 | 0 | Factual
increased total bilirubin | 0 | 0 | Factual
increased direct bilirubin | 0 | 0 | Factual
increased AST | 0 | 0 | Factual
increased ALT | 0 | 0 | Factual
increased PSA | 0 | 0 | Factual
increased white blood cell count | 0 | 0 | Factual
no hydronephrosis | 0 | 0 | Factual
empty bladder | 0 | 0 | Factual
traces of blood in bladder catheter | 0 | 0 | Factual
no urologic surgery | 0 | 0 | Negated
prostatic hypertrophy | -672 | 0 | Factual
overactive bladder | -672 | 0 | Factual
recurrent prostatitis | -672 | 0 | Factual
use of statins | 0 | 0 | Negated
volume expansion | 0 | 504 | Factual
diuretic treatment | 0 | 504 | Factual
alpha-agonist | 0 | 504 | Factual
antibiotic treatment | 0 | 504 | Factual
furosemide | 0 | 192 | Factual
femoral central venous catheter | 0 | 0 | Factual
HFR-Supra | 0 | 120 | Factual
endogenous reinfusion | 0 | 120 | Factual
myoglobin removal | 0 | 120 | Factual
inflammatory status reduction | 0 | 120 | Factual
fluid balance maintenance | 0 | 120 | Factual
ultrafiltration | 0 | 120 | Factual
adsorbent cartridge | 0 | 120 | Factual
low molecular weight heparin | 0 | 0 | Factual
myoglobin reduction | 0 | 120 | Factual
CPK reduction | 0 | 120 | Factual
LDH reduction | 0 | 120 | Factual
CRP reduction | 0 | 120 | Factual
PCT reduction | 0 | 120 | Factual
urine output increase | 96 | 192 | Factual
furosemide tapering | 192 | 192 | Factual
antibiotic therapy change | 0 | 504 | Factual
piperacillin/tazobactam | 0 | 120 | Factual
meropenem | 120 | 504 | Factual
femoral hemodialysis catheter removal | 120 | 120 | Factual
right jugular central venous catheter placement | 120 | 120 | Factual
on-line hemodiafiltration | 120 | 168 | Factual
high-flux hemodialysis | 168 | 192 | Factual
dialysis discontinuation | 504 | 504 | Factual
urea reduction | 504 | 504 | Factual
creatinine reduction | 504 | 504 | Factual
CRP reduction | 504 | 504 | Factual
total bilirubin reduction | 504 | 504 | Factual
ASL reduction | 504 | 504 | Factual
ALT reduction | 504 | 504 | Factual
PSA reduction | 504 | 504 | Factual
white blood cell count reduction | 504 | 504 | Factual
hospital discharge | 504 | 504 | Factual
urea follow-up | 1008 | 1008 | Factual
creatinine follow-up | 1008 | 1008 | Factual
GFR follow-up | 1008 | 1008 | Factual