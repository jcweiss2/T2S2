56 years old | 0
woman | 0
admitted to the hospital | -1440
schizophrenia | -1440
perforated diverticulitis | -1440
sigmoid resection | -1440
anastomotic leak | -1440
defunctioning ileostomy | -1440
feculent peritonitis | -1440
surgical wound dehiscence | -1440
percutaneous drainage | -1440
laparotomy | -1440
prolonged broad-spectrum antibiotic treatment | -1440
wound debridements | -1440
high-protein/caloric diet | -1440
poor oral intake | -1440
acetaminophen 650 mg 4 times per day | -1440
acetaminophen dose increased to 650 mg every 4 hours | -1440
hypovolemic shock | -1440
high gastrointestinal losses | -1440
transferred to intensive care unit | 0
new abdominal collections | 0
acute kidney injury (AKI) | 0
high-anion-gap metabolic acidosis (HAGMA) | 0
negative alcohol screen | 0
normal liver function tests | 0
lactate | 0
negative salicylates | 0
mildly elevated beta-hydroxybutyrate | 0
elevated anion gap | 0
elevated serum osmolal gap | 0
acetaminophen stopped | 0
volume expansion with dextrose and bicarbonate drip | 0
N-acetyl cysteine administered | 0
sustained low-efficiency dialysis (SLED) initiated | 0
markedly increased excretion of 5-oxoproline | 24
HAGMA improved | 24
continued vasopressor support | 48
continued ventilatory support | 48
ventilator-associated pneumonia | 48
transferred back to medical ward | 48
recurrent aspirations | 72
passed away | 72
