57 years old | 0
female | 0
family history of mitral valve prolapse | 0
admitted to the hospital | 0
altered mental status | 0
fatigue | -168
generalized weakness | -168
nonbloody vomiting | -168
diarrhea | -168
denies chest pressure | 0
denies chest pain | 0
denies fever | 0
denies history of intravenous drug use | 0
heart rate of 135 beats per minute | 0
Janeway lesions | 0
Osler nodes | 0
splinter hemorrhages | 0
white blood cell count of 17 000/mm3 | 0
hemoglobin of 11.7 g/dL | 0
platelets 89 000/mm3 | 0
point of care troponin of 0.28 ng/mL | 0
sinus tachycardia | 0
nonspecific ST-wave changes | 0
blood cultures drawn | 0
intravenous fluids | 0
empiric intravenous antibiotics | 0
ceftriaxone | 0
vancomycin | 0
follow-up troponin of 0.85 | 12
heparin drip | 12
chest pain free | 12
persistent sinus tachycardia | 12
no ST-segment changes | 12
subacute infarcts in the cerebral hemispheres | 12
infarctions in the kidney and spleen | 12
heparin drip stopped | 12
transthoracic echocardiogram | 12
cardiology consulted | 12
blood cultures positive for methicillin-sensitive Staphylococcus aureus | 24
ejection fraction of 55% | 24
no vegetations | 24
chest pain | 48
new diffuse ST-segment elevation | 48
PR depression | 48
pericarditis | 48
nonsteroidal anti-inflammatory drugs | 48
repeat TTE | 48
ejection fraction of 35% to 40% | 48
severe diffuse hypokinesis of the apical wall | 48
possible vegetation on mitral valve | 48
transesophageal echocardiogram | 72
ejection fraction of 30% to 35% | 72
severe hypokinesis | 72
medium-sized vegetation on the atrial aspect of the tip of the anterior leaflet of mitral valve | 72
moderate to severe mitral valve regurgitation | 72
cardiothoracic surgery consulted | 72
shortness of breath | 72
cardiogenic shock | 72
vasopressor support | 72
troponin of 49.50 ng/mL | 72
emergent cardiac catheterization | 72
100% occlusion of the proximal left anterior descending artery | 72
septic embolus | 72
mitral valve replacement | 96
coronary artery bypass grafting | 96
gross specimen showed vegetations involving the mitral valve leaflets | 96
discharged to a rehabilitation center | 336
intravenous antibiotics | 336
metoprolol tartrate | 336
furosemide | 336
potassium chloride | 336
seizure | 504
pulseless electrical activity | 504
cardiopulmonary resuscitation | 504
return of spontaneous circulation | 504
potassium of 8 | 504
elevated troponins | 504
lactic acid | 504
evolution of the previously known ischemic infarctions | 504
no acute or hemorrhagic components | 504
stat TTE postcardiac arrest | 504
ejection fraction of 20% | 504
cardiac arrest likely secondary to seizure | 504
hyperkalemia | 504
terminally extubated | 510