40 years old | 0
female | 0
chronic alcoholic | 0
admitted to the hospital | 0
found sleeping in a car on the street | -1
drinking alcohol on a daily basis | -24
last drink was 1 h prior to arrival | -1
hypothermic at 81°F on arrival | 0
warming blanket | 0
improved to 91.7°F | 1
improved to 97°F | 8
white blood cell count of 9.1 | 0
mild left shift | 0
hemoglobin 11 | 0
hematocrit 34 | 0
platelets 458 | 0
serum alcohol level 0.01 | 0
creatinine phosphokinase 564 | 0
blood urea nitrogen 16 | 0
creatinine 0.4 | 0
glucose 58 | 0
aspartate transaminase 188 | 0
alanine transaminase 69 | 0
alkaline phosphatase 216 | 0
TSH 1.07 | 0
prolactin 44.9 | 0
amylase 498 | 0
lipase 1,200 | 0
ammonia 26 | 0
serum carboxyhemoglobin level 2.4 | 0
magnesium 1.3 | 0
cortisol 38 | 0
β-HCG negative | 0
witnessed generalized tonic-clonic seizure | 2
intravenous lorazepam 2 mg | 2
loading dose of levetiracetam 1,000 mg | 2
transient hypotension | 2
fluid challenge | 2
normal saline | 2
vancomycin | 2
cefepime | 2
metronidazole | 2
sepsis workup | 4
antibiotics held off | 4
sonogram (abdomen) | 4
fatty liver | 4
trace ascites | 4
CAT scan (abdomen and pelvis) | 8
peripancreatic fluid | 8
fluid in the splenic flexure of the colon | 8
fluid in the inferior aspect of the spleen | 8
pancreas symmetrically enhanced | 8
no evidence of pancreatic necrosis | 8
no evidence of hemorrhage | 8
no evidence of peripancreatic abscess | 8
no evidence of pancreatic mass | 8
medically managed | 12
discharged from hospital | 96
low-fiber low-fat diet | 96