74 years old | 0  
    male | 0  
    presented with a one-month history of worsening pruritus | -720  
    confusion | -720  
    multiple falls | -720  
    fever | -720  
    lethargy | -720  
    night sweats | -720  
    previous coronary stenting for ischaemic heart disease | 0  
    taking aspirin | 0  
    non-smoker | 0  
    occasionally consumed alcohol | 0  
    pyrexial | 0  
    tachycardic | 0  
    deranged liver function | 0  
    bilirubin 28 | 0  
    alanine transaminase 106 | 0  
    alkaline phosphatase 600 | 0  
    synthetic impairment | 0  
    INR 2.0 | 0  
    albumin 29 | 0  
    pancytopenia | 0  
    hemoglobin 85 | 0  
    white cell count 2.7 | 0  
    platelets 71 | 0  
    raised C-reactive protein 55 | 0  
    initiated on co-amoxiclav for biliary sepsis | 0  
    abdominal ultrasound showed thickened gallbladder without stones | 0  
    no biliary duct dilatation | 0  
    normal liver | 0  
    portal venous flow | 0  
    spleen enlarged at 16 cm | 0  
    hypoechoic area 30x43 mm | 0  
    CT abdomen confirmed enlarged spleen | 0  
    magnetic resonance cholangiopancreatography normal | 0  
    work-up for acute liver injury | 0  
    viral serology | 0  
    autoimmune screen | 0  
    immunoglobulins | 0  
    blood cultures negative | 0  
    continued to spike fevers | 96  
    haemodynamic instability | 96  
    two medical emergency calls | 96  
    antibiotics escalated to piperacillin/tazobactam | 96  
    raised lactate | 96  
    worsening pancytopenia | 96  
    acute kidney injury | 96  
    deterioration in liver function | 96  
    jaundice | 96  
    INR up to 2.0 | 96  
    lactate dehydrogenase >2000 IU/L | 96  
    ferritin >3000 ug/L | 96  
    staging CT showed bilateral pleural effusions | 96  
    minimal ascites | 96  
    peri-pancreatic stranding suggestive of mild pancreatitis | 96  
    amylase marginally raised at 125 iu/L | 96  
    bone marrow aspirate | 96  
    trephine biopsy | 96  
    development of hepatic encephalopathy | 96  
    hypoxia | 96  
    hypotensive | 96  
    persistent tachycardia | 96  
    fluid resuscitation | 96  
    antibiotics escalated to meropenem | 96  
    hepatology review recommended viral serology tests | 96  
    hepatitis A negative | 96  
    hepatitis E negative | 96  
    hepatitis B core antibody negative | 96  
    leptospirosis negative | 96  
    brucella negative | 96  
    herpes simplex virus serology negative | 96  
    preliminary bone marrow biopsy showed reactive changes | 96  
    no evidence of lymphoma | 96  
    no haemophagocytosis | 96  
    deterioration with multi-organ failure | 264  
    clinical diagnosis of haemophagocytic lymphohistiocytosis | 264  
    met HLH-2004 criteria | 264  
    splenomegaly | 264  
    fever >38.5 | 264  
    cytopenia | 264  
    hemoglobin <90 g/l | 264  
    platelets <100×10^9/l | 264  
    hypertriglyceridemia ≥3.0 mmol/l | 264  
    ferritin >500 ng/ml | 264  
    administration of 1g methylprednisolone | 264  
    rapid deterioration | 264  
    pH 6.89 | 264  
    lactate 17.8 | 264  
    consensus of imminent death | 264  
    passed away | 264  
    bone marrow trephine biopsy confirmed diffuse large B-cell lymphoma | 264  
    80% blast | 264  
    confirming haemophagocytic lymphohistiocytosis with underlying malignancy | 264  
    patient died | 264  