55 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
morbidly obese | 0 | 0 | Factual
diabetes mellitus | 0 | 0 | Factual
end-stage renal disease | 0 | 0 | Factual
hemodialysis | 0 | 0 | Factual
peripheral vascular disease | 0 | 0 | Factual
left below knee amputation | 0 | 0 | Factual
right above knee amputation | 0 | 0 | Factual
right extra anatomical axillobifemoral bypass graft | 0 | 0 | Factual
admitted to emergency department | 0 | 0 | Factual
right-sided abdominal pain | -48 | 0 | Factual
vomiting | -48 | 0 | Factual
fever | -48 | 0 | Factual
conscious | 0 | 0 | Factual
alert | 0 | 0 | Factual
oriented | 0 | 0 | Factual
pale | 0 | 0 | Factual
sick | 0 | 0 | Factual
temperature 37.8°C | 0 | 0 | Factual
blood pressure 150/90 mmHg | 0 | 0 | Factual
oxygen saturation 95% | 0 | 0 | Factual
abdomen distended | 0 | 0 | Factual
tympanic | 0 | 0 | Factual
right upper quadrant tenderness | 0 | 0 | Factual
right flank tenderness | 0 | 0 | Factual
total leukocyte count 20 × 10^3 | 0 | 0 | Factual
hemoglobin 10.7 gm% | 0 | 0 | Factual
acidotic pH 7.33 | 0 | 0 | Factual
laboratory evidence of end-stage renal disease | 0 | 0 | Factual
air under the right hemi-diaphragm | 0 | 0 | Factual
perforated viscous | 0 | 0 | Possible
computed tomography scan | 0 | 0 | Factual
right perinephric collection | 0 | 0 | Factual
extension into the right sub-phrenic region | 0 | 0 | Factual
gas in the right collecting system | 0 | 0 | Factual
gas in the urinary bladder | 0 | 0 | Factual
no gas in the renal parenchyma | 0 | 0 | Factual
right atrial thrombus | 0 | 0 | Factual
parenteral antibiotics | 0 | 0 | Factual
admitted to intensive care unit | 0 | 0 | Factual
percutaneous drainage | 0 | 0 | Factual
failed percutaneous drainage | 0 | 0 | Factual
not fit for general anesthesia | 0 | 0 | Factual
open drainage | 0 | 0 | Factual
loculated perinephric and sub-phrenic collection | 0 | 0 | Factual
cystoscopy | 0 | 0 | Factual
abnormal bladder mucosa | 0 | 0 | Factual
multiple cystic lesions | 0 | 0 | Factual
air “bubbles” in the bladder | 0 | 0 | Factual
ureteric Double J stent | 0 | 0 | Factual
urethral catheter | 0 | 0 | Factual
reasonably well during the procedure | 0 | 0 | Factual
condition deteriorated | 24 | 48 | Factual
culture of the collection | 24 | 48 | Factual
Klebsiella pneumonia extended-spectrum β-lactamase | 24 | 48 | Factual
severe sepsis | 48 | 48 | Factual
multiple organ failure | 48 | 48 | Factual
died | 48 | 48 | Factual