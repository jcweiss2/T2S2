5 years old | 0
female | 0
admitted to the pediatric intensive care unit | 0
cough | -336
fever | -120
headache | -24
vomiting | -24
altered interactions | -24
retarded height growth | -8760
decreased activity | -8760
uncomplicated birth | -43800
normal growth | -43800
temperature of 38.7°C | 0
heart rate of 105 beats per minute | 0
respiratory rate of 35 breaths per minute | 0
blood pressure of 90/55 mmHg | 0
oxyhemoglobin saturation of 90% | 0
generalized puffiness | 0
non-pitting edema | 0
capillary refilled time >3 seconds | 0
rales | 0
normal cardiac auscultation | 0
soft abdomen | 0
mildly distended abdomen | 0
normal bowel sounds | 0
slightly confused | 0
could not properly respond to commands | 0
hemoglobin level of 97 g/L | 0
white blood cell count of 2.5×10^9/L | 0
neutrophils 70% | 0
blood platelet 75×10^9/L | 0
normal electrolytes | 0
normal glucose | 0
normal albumin | 0
normal creatine kinase | 0
normal blood gas | 0
left lobe pneumonia | 0
mild pleural effusion | 0
mild pericardial effusion | 0
normal cardiac ejection fraction | 0
normal MRI scan of the brain | 0
normal cerebrospinal fluid exam | 0
diagnosed as pneumonia | 0
diagnosed as sepsis | 0
empiric antibiotic therapy | 0
immunoglobulin supply | 0
restricted fluid administration | 0
comatose | 24
temperature dropped to 35°C | 24
hypotension | 24
arrhythmia | 24
hypoxia | 24
SaO2 decreased to 75% | 24
prolonged Q–T interval | 24
thyroid studies ordered | 0
thyroxin undetectable | 24
TSH extremely high | 24
elevated anti-thyroid peroxidase | 48
elevated anti-thyroglobulin | 48
mild bilateral thyroid enlargement | 48
small tubercles in the left thyroid | 48
diagnosed with myxedema coma | 24
hormone replacement started | 24
intravenous dexamethasone | 24
oral levothyroxine | 24
vasopressor | 24
mechanical ventilation | 24
continuous renal replacement treatment | 24
consciousness restored | 48
temperature returned to normal | 48
extubated | 120
dosage of oral levothyroxine reduced | 336
discharged | 336
height increased 9 cm | 4032
more active | 4032
father diagnosed with Hashimoto's thyroiditis | 4032
grandmother diagnosed with Hashimoto's thyroiditis | 4032