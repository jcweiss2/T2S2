76 years old | 0
male | 0
admitted to the Emergency Department | 0
psoriasis | -6720
chronic kidney disease stage 4 | -6720
essential hypertension | -6720
amlodipine | -6720
atenolol | -6720
lowered level of awareness | 0
sustained bradycardia | 0
denied syncope | 0
denied angina | 0
denied palpitation | 0
heart rate of 26 beats per minute | 0
blood pressure of 80/40 mmHg | 0
mean arterial pressure of 53 mmHg | 0
body temperature of 35.6°C | 0
respiratory rate of 18 breaths per minute | 0
peripheral oxygen saturation of 95% | 0
white blood cell count of 5.450 cells/μL | 0
creatinine level of 3.7 mg/dL | 0
serum potassium level of 7.3 mg/dL | 0
TSH of 4.92 μUI/mL | 0
C-reactive protein of 48.9 mg/dL | 0
normal chest X-ray | 0
normal systolic and diastolic function | 0
no remarkable changes with the heart valves | 0
sinus bradycardia with junctional escape rhythm | 0
hypothesis of BRASH syndrome | 0
intravenous bolus of sodium chloride | 0
atropine | 0
glucagon | 0
calcium gluconate | 0
hydrocortisone | 0
sodium bicarbonate | 0
dextrose with insulin | 0
suspension of previous medications | 0
continuous infusion of epinephrine | 0
temporary transvenous pacemaker | 24
admitted to the Intensive Care Unit | 0
correction of hyperkalemia | 24
return of creatinine levels to baseline values | 96
suspension of epinephrine infusion | 96
removal of temporary pacemaker | 120
discharged | 192
normal sinus rhythm | 192
serum creatinine of 2.36 mg/dL | 192
potassium of 4.9 mg/dL | 192