39 years old | 0
female | 0
32 weeks of gestation | 0
admitted to the emergency room | 0
shortness of breath | 0
progressive limb weakness | 0
2-year history of worsening neck pain | -8760
weakness in her right arm | -120
weakness in her left arm | -60
weakness in both legs | -60
numbness from the neck down | -60
fever | -72
no complaints of anosmia | 0
no complaints of seizure | 0
no complaints of blurred vision | 0
no complaints of slurred speech | 0
no complaints of dysphagia | 0
no complaints of hoarseness | 0
no complaints of skewed face | 0
no urination or defecation disturbances | 0
history of contraceptive injection for 15 years | -13140
consumed ibuprofen and paracetamol for neck pain for 2 years | -8760
intact mental status | 0
no meningeal signs | 0
no cranial nerve palsy | 0
tetraplegia | 0
hypoesthesia below the C3–C4 spinal cord segments | 0
abnormal proprioception | 0
increased tendon reflexes | 0
positive Babinski and Chaddock reflexes | 0
PCR testing of a nasopharyngeal swab was positive for COVID-19 | 0
chest radiography revealed paracardial infiltrates | 0
respiratory failure | 0
increased D-dimer | 0
hypokalemia | 0
admitted to the intensive care unit | 0
intubated | 0
treated with high-dose n-acetylcysteine | 0
treated with remdesivir | 0
treated with zinc | 0
treated with vitamin D | 0
treated with vitamin C | 0
emergency cesarean section | 24
tumor excision by craniotomy | 48
histopathological examination revealed transitional and angiomatous type WHO grade 1 meningioma | 48
patient's awareness increased briefly after surgery | 48
patient's condition continued to deteriorate | 72
blood pressure decreased to 60/30 mmHg | 72
administered norepinephrine | 72
septic shock | 96
respiratory failure | 96
patient died | 120