74 years old | 0
male | 0
admitted to the hospital | 0
pruritus | -720
confusion | -720
multiple falls | -720
fever | -720
lethargy | -720
night sweats | -720
ischaemic heart disease | -720
coronary stenting | -720
aspirin | -720
non-smoker | 0
occasionally consumed alcohol | 0
pyrexial | 0
tachycardic | 0
abdominal examination unremarkable | 0
deranged liver function | 0
Bilirubin 28 | 0
Alanine transaminase 106 | 0
Alkaline phosphatase 600 | 0
synthetic impairment | 0
INR 2.0 | 0
Albumin 29 | 0
pancytopenia | 0
Haemoglobin 85 | 0
White Cell Count 2.7 | 0
Platelets 71 | 0
C-reactive protein 55 | 0
co-amoxiclav | 0
biliary sepsis | 0
abdominal ultrasound | 0
thickened gallbladder | 0
no stones | 0
no biliary duct dilatation | 0
normal liver | 0
normal portal venous flow | 0
enlarged spleen | 0
hypoechoic area | 0
CT abdomen | 0
magnetic resonance cholangiopancreatography | 0
normal | 0
viral serology | 0
autoimmune screen | 0
immunoglobulins | 0
unrevealing | 0
blood cultures | 0
negative | 0
spiking temperature | 0
Piperacillin/Tazobactam | 96
haemodynamic instability | 96
medical emergency calls | 96
raised lactate | 96
worsening pancytopenia | 96
acute kidney injury | 96
deterioration in liver function | 96
jaundice | 96
INR up to 2.0 | 96
Lactate dehydrogenase >2000 IU/L | 96
ferritin >3000 ug/L | 96
staging CT | 96
new bilateral pleural effusions | 96
minimal ascites | 96
peri-pancreatic stranding | 96
mild pancreatitis | 96
amylase 125 iu/L | 96
bone marrow aspirate | 96
trephine biopsy | 96
hepatic encephalopathy | 120
hypoxia | 120
hypotensive | 120
persistent tachycardia | 120
fluid resuscitation | 120
Meropenem | 120
hepatology review | 120
Hepatitis A | 120
Hepatitis E | 120
Hepatitis B core antibody | 120
leptospirosis | 120
Brucella | 120
herpes simplex virus serology | 120
normal | 120
preliminary bone marrow biopsy results | 120
reactive changes | 120
infection | 120
no evidence of lymphoma | 120
no haemophagocytosis | 120
clinical diagnosis of haemophagocytic lymphohistiocytosis | 264
methylprednisolone | 264
family’s consent | 264
deteriorated rapidly | 264
imminent death | 264
pH 6.89 | 264
Lactate 17.8 | 264
passed away | 264
bone marrow trephine biopsy result | 264
diffuse large B-cell lymphoma | 264
80% blast | 264
haemophagocytic lymphohistiocytosis | 264
underlying malignancy | 264