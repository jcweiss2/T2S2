77 years old | 0
    female | 0
    admitted to ICU | 0
    bilateral pneumonia | 0
    acute kidney injury | 0
    intubated | 0
    respiratory distress | 0
    subclavian central line inserted | 0
    vasopressors started | 0
    piperacillin/tazobactam initiated | 0
    clindamycin initiated | 0
    meropenem initiated | -96
    teicoplanin initiated | -96
    rising leukocyte counts | -96
    colistin initiated | -168
    carbapenem resistant organism in endotracheal secretions | -168
    fluconazole initiated | -120
    watery diarrhea | -144
    racecadotril initiated | -144
    metronidazole initiated | -144
    Saccharomyces sachet initiated | -144
    antibiotic-induced diarrhea suspected | -144
    Clostridium difficile infection suspected | -144
    stool routine/microscopy negative | -144
    stool culture negative | -144
    C. difficile toxin negative | -144
    diarrhea resolved | -144
    hypotension | -168
    diarrhea recurrence | -168
    caspofungin initiated | -168
    fluconazole discontinued | -168
    cultures repeated | -168
    blood culture sterile (48 hours) | -144
    Saccharomyces cerevisiae in central line blood | -192
    Saccharomyces cerevisiae in peripheral blood | -192
    caspofungin discontinued | -192
    amphotericin B initiated | -192
    Saccharomyces sachet discontinued | -192
    central line removed | -192
    repeat blood cultures negative (3rd day) | -216
    repeat blood cultures negative (7th day) | -288
    death | 576
    uncontrolled diabetes (HbA1c 8.4) | 0
    hypertension | 0
    chronic obstructive airway disease | 0
    no fungal growth in repeat cultures | -216
    no fungal growth in repeat cultures | -288
    mechanical ventilation | 0
    probiotic contamination risk | 0
    immune compromised status | 0
    broad-spectrum antibiotics use | 0
    invasive lines | 0
    long hospital stay | 0
    probiotics discontinued | -192
    antifungal treatment | -192
    catheter tip culture recommended | 0
    clinician awareness required | 0
    MIC breakpoint undefined | 0
    echinocandin studies needed | 0
    warning tags for manufacturers | 0
    differentiation from Candida required | 0
    Lactobacillus probiotics preferred | 0
    Saccharomyces fungemia risk factors | 0
    antifungal susceptibility tested | -192
    amphotericin B effective | -192
    patient on Saccharomyces supplements | -144
    probiotics used in ICU | 0
    critical illness | 0
    fungemia | -192
    septic shock | -192
    invasive fungal infection | -192
    antifungal therapy adjustment | -192
    line removal for infection control | -192
    hypotension management | -168
    diarrhea management | -144
    antifungal switch | -168
    stool testing performed | -144
    blood cultures sent | -144
    probiotic administration | -144
    risk factor assessment | 0
    mortality | 576
    no evidence of C. difficile | -144
    negative stool studies | -144
    positive blood cultures | -192
    yeast identification | -192
    treatment discontinuation | -192
    line removal | -192
    antifungal efficacy | -192
    negative follow-up cultures | -216
    negative follow-up cultures | -288
    death after 24 days | 576
    probiotic-related complications | -192
    fungemia source investigation | -192
    literature review | -192
    antifungal choice dilemma | -192
    MIC breakpoint uncertainty | 0
    amphotericin B selection | -192
    probiotics handling precautions | 0
    Saccharomyces risk awareness | 0
    Lactobacillus alternative | 0
    central line colonization risk | 0
    gut translocation risk | 0
    ICU precautions | 0
    patient monitoring | 0
    infection control measures | -192
    antifungal combination use | 0
    mortality risk factors | 0
    no Candida differentiation | 0
    antifungal susceptibility report available | -192
    Saccharomyces confirmed | -192
    probiotics stopped | -192
    invasive procedures | 0
    immunocompromised state | 0
    uncontrolled diabetes as risk | 0
    chronic lung disease | 0
    mechanical ventilation as risk | 0
    broad-spectrum antibiotics as risk | 0
    line removal for fungemia | -192
    antifungal therapy change | -168
    negative blood cultures initially | -144
    positive blood cultures later | -192
    yeast growth identification | -192
    antifungal adjustment | -192
    line removal confirmation | -192
    probiotics cessation | -192
    amphotericin B effectiveness | -192
    follow-up cultures | -216
    follow-up cultures | -288
    patient outcome | 576
    probiotic-induced fungemia | -192
    line-related infection | -192
    gut translocation hypothesis | -192
    risk factor mitigation | 0
    treatment protocol adherence | 0
    mortality despite treatment | 576
    no further fungal growth post-treatment | -216
    no further fungal growth post-treatment | -288
    death after prolonged ICU stay | 576
    antifungal therapy initiated | -120
    antifungal therapy adjustment | -168
    antifungal therapy change to amphotericin | -192
    treatment discontinuation | -192
    probiotic administration complications | -144
    Saccharomyces fungemia diagnosis | -192
    line removal as intervention | -192
    amphotericin B as treatment | -192
    negative follow-up cultures | -216
    negative follow-up cultures | -288
    death due to complications | 576
    uncontrolled diabetes management | 0
    hypertension management | 0
    chronic obstructive airway disease management | 0
    bilateral pneumonia management | 0
    acute kidney injury management | 0
    respiratory distress management | 0
    vasopressor management | 0
    antibiotic therapy adjustments | -96
    antibiotic therapy adjustments | -168
    antifungal therapy adjustments | -120
    antifungal therapy adjustments | -168
    probiotic administration | -144
    diarrhea treatment | -144
    hypotension treatment | -168
    line removal procedure | -192
    infection source control | -192
    antifungal selection | -192
    patient monitoring post-intervention | -216
    patient monitoring post-intervention | -288
    mortality documentation | 576
    no evidence of C. difficile infection | -144
    stool studies negative | -144
    blood culture positivity | -192
    yeast species identification | -192
    treatment alteration | -192
    line removal confirmation | -192
    amphotericin B efficacy | -192
    follow-up culture negativity | -216
    follow-up culture negativity | -288
    death after 24 days | 576
    probiotic cessation | -192
    line removal success | -192
    amphotericin B administration | -192
    negative repeat cultures | -216
    negative repeat cultures | -288
    mortality despite interventions | 576
    Saccharomyces fungemia confirmation | -192
    risk factor presence | 0
    appropriate antifungal use | -192
    infection control measures | -192
    treatment adherence | 0
    patient outcome monitoring | 0
    death confirmation | 576
    no further complications post-treatment | -216
    no further complications post-treatment | -288
    antifungal therapy success | -216
    antifungal therapy success | -288
    mortality despite antifungal therapy | 576
    probiotic-related fungemia | -192
    line-related fungemia | -192
    gut translocation possibility | -192
    risk factor documentation | 0
    treatment protocol followed | 0
    death due to fungemia | 576
    prolonged ICU stay | 576
    no improvement post-treatment | 576
    death after interventions | 576
    Saccharomyces fungemia as cause | -192
    risk factors contributing | 0
    appropriate management steps | -192
    line removal contributing | -192
    amphotericin B as appropriate | -192
    negative follow-up cultures indicating control | -216
    negative follow-up cultures indicating control | -288
    death despite control measures | 576
    probiotic discontinuation effect | -192
    line removal effect | -192
    antifungal therapy effect | -192
    mortality risk factors | 0
    uncontrolled diabetes contributing | 0
    chronic lung disease contributing | 0
    mechanical ventilation contributing | 0
    broad-spectrum antibiotics contributing | 0
    invasive lines contributing | 0
    long ICU stay contributing | 0
    immunocompromised state contributing | 0
    Saccharomyces fungemia complications | -192
    septic shock contributing | -192
    hypotension contributing | -168
    diarrhea contributing | -144
    fungemia contributing | -192
    amphotericin B administration | -192
    caspofungin discontinuation | -192
    fluconazole discontinuation | -168
    probiotic cessation | -192
    central line removal | -192
    negative follow-up cultures | -216
    negative follow-up cultures | -288
    death outcome | 576
    no Candida differentiation | 0
    Saccharomyces identification | -192
    antifungal susceptibility testing | -192
    MIC breakpoint undefined | 0
    echinocandin studies needed | 0
    warning tags for probiotics | 0
    Lactobacillus preference | 0
    clinician awareness | 0
    catheter tip culture recommendation | 0
    manufacturer warnings | 0
    MIC definition needed | 0
    echinocandin research needed | 0
    probiotic handling precautions | 0
    risk factor awareness | 0
    differentiation from Candida importance | 0
    treatment strategy adherence | 0
    mortality documentation | 576
    death after 24 days | 576
    no survival post-treatment | 576
    antifungal therapy failure | 576
    fungemia persistence | -192
    septic shock persistence | -192
    hypotension persistence | -168
    diarrhea recurrence persistence | -168
    Saccharomyces persistence | -192
    amphotericin B administration | -192
    line removal persistence | -192
    probiotic discontinuation persistence | -192
    negative cultures post-treatment | -216
    negative cultures post-treatment | -288
    death despite negative cultures | 576
    prolonged ICU stay contributing | 576
    risk factor accumulation | 0
    uncontrolled diabetes as risk | 0
    chronic lung disease as risk | 0
    mechanical ventilation as risk | 0
    invasive lines as risk | 0
    broad-spectrum antibiotics as risk | 0
    immunocompromised state as risk | 0
    Saccharomyces fungemia confirmation | -192
    amphotericin B administration | -192
    line removal confirmation | -192
    probiotic discontinuation confirmation | -192
    negative follow-up cultures confirmation | -216
    negative follow-up cultures confirmation | -288
    death confirmation | 576
    no further intervention impact | 576
    mortality final | 576
    death due to complications | 576
    fungemia as primary cause | -192
    risk factors contributing | 0
    management steps taken | -192
    no survival | 576
    death after 24 days | 576
    ICU mortality | 576
    fungemia-related death | 576
    probiotic-related death | 576
    Saccharomyces complications | -192
    risk factor presence | 0
    treatment adherence | 0
    line removal adherence | -192
    antifungal adherence | -192
    probiotic discontinuation adherence | -192
    negative cultures post-treatment | -216
    negative cultures post-treatment | -288
    death outcome final | 576
    death after interventions | 576
    no improvement | 576
    mortality documentation final | 576
    death after 24 days | 576
    ICU stay duration | 576
    prolonged hospitalization | 576
    death despite treatment | 576
    fungemia as mortality cause | -192
    risk factors contributing | 0
    management steps insufficient | 576
    death inevitable | 576
    no recovery | 576
    patient demise | 576
    death after prolonged stay | 576
    ICU complications | 576
    fungemia complications | 576
    septic shock complications | 576
    hypotension complications | 576
    diarrhea complications | 576
    Saccharomyces complications | 576
    amphotericin B administration insufficient | 576
    line removal insufficient | 576
    probiotic discontinuation insufficient | 576
    negative cultures insufficient | 576
    death despite negative cultures | 576
    mortality documentation | 576
    death after 24 days | 576
    ICU mortality | 576
    fungemia-related mortality | 576
    probiotic-related mortality | 576
    risk factor-related mortality | 0
    uncontrolled diabetes mortality impact | 0
    chronic lung disease mortality impact | 0
    mechanical ventilation mortality impact | 0
    invasive lines mortality impact | 0
    broad-spectrum antibiotics mortality impact | 0
    immunocompromised state mortality impact | 0
    Saccharomyces mortality impact | -192
    amphotericin B impact | -192
    line removal impact | -192
    probiotic discontinuation impact | -192
    negative cultures impact | -216
    negative cultures impact | -288
    death despite interventions | 576
    mortality final | 576
    death after 24 days | 576
    ICU stay end | 576
    patient outcome final | 576
    death documentation | 576
    no survival post-ICU | 576
    death confirmed | 576
    mortality conclusion | 576
    death due to fungemia | 576
    risk factors conclusion | 0
    management steps conclusion | 0
    antifungal therapy conclusion | 0
    line removal conclusion | 0
    probiotic discontinuation conclusion | 0
    negative cultures conclusion | 0
    death conclusion | 576
    Saccharomyces fungemia conclusion | -192
    ICU mortality conclusion | 576
    probiotic-related death conclusion | 576
    risk factor accumulation conclusion | 0
    uncontrolled diabetes conclusion | 0
    chronic lung disease conclusion |4
    0
    chronic obstructive airway disease | 0
    hypertension | 0
    bilateral pneumonia | 0
    acute kidney injury | 0
    intubation | 0
    respiratory distress | 0
    subclavian central line insertion | 0
    vasopressors initiation | 0
    piperacillin/tazobactam initiation | 0
    clindamycin initiation | 0
    meropenem initiation | -96
    teicoplanin initiation | -96
    leukocyte count elevation | -96
    colistin initiation | -168
    carbapenem resistant organism detection | -168
    fluconazole initiation | -120
    diarrhea onset | -144
    racecadotril initiation | -144
    metronidazole initiation | -144
    Saccharomyces sachet initiation | -144
    antibiotic-associated diarrhea suspicion | -144
    Clostridium difficile suspicion | -144
    stool tests negative | -144
    diarrhea resolution | -144
    hypotension onset | -168
    diarrhea recurrence | -168
    caspofungin initiation | -168
    fluconazole discontinuation | -168
    repeat cultures | -168
    sterile blood cultures (48 hours) | -144
    Saccharomyces cerevisiae in central line blood | -192
    Saccharomyces cerevisiae in peripheral blood | -192
    caspofungin discontinuation | -192
    amphotericin B initiation | -192
    Saccharomyces sachet discontinuation | -192
    central line removal | -192
    repeat blood cultures negative (3rd day) | -216
    repeat blood cultures negative (7th day) | -288
    death | 576
    uncontrolled diabetes (HbA1c 8.4) | 0
    hypertension | 0
    chronic obstructive airway disease | 0
    mechanical ventilation | 0
    immune compromised status | 0
    invasive lines | 0
    broad-spectrum antibiotic use | 0
    long hospital stay | 0
    probiotic contamination risk | 0
    probiotics discontinued | -192
    antifungal treatment initiation | -192
    catheter tip culture recommendation | 0
    clinician awareness needed | 0
    MIC breakpoint undefined | 0
    echinocandin studies needed | 0
    warning tags for manufacturers | 0
    differentiation from Candida | 0
    Lactobacillus preference | 0
    Saccharomyces fungemia risk factors | 0
    antifungal susceptibility tested | -192
    amphotericin B effectiveness | -192
    probiotics used in ICU | 0
    critical illness | 0
    fungemia | -192
    septic shock | -192
    invasive fungal infection | -192
    antifungal therapy adjustment | -192
    line removal for infection control | -192
    hypotension management | -168
    diarrhea management | -144
    antifungal switch | -168
    stool testing performed | -144
    blood cultures sent | -144
    probiotic administration | -144
    risk factor assessment | 0
    mortality | 576
    no C. difficile infection | -144
    negative stool studies | -144
    positive blood cultures | -192
    yeast identification | -192
    treatment discontinuation | -192
    line removal | -192
    antifungal efficacy | -192
    negative follow-up cultures | -216
    negative follow-up cultures | -288
    death after 24 days | 576
    probiotic-related complications | -192
    fungemia source investigation | -192
    literature review | -192
    antifungal choice dilemma | -192
    MIC breakpoint uncertainty | 0
    amphotericin B selection | -192
    probiotics handling precautions | 0
    Saccharomyces risk awareness | 0
    Lactobacillus alternative | 0
    central line colonization risk | 0
    gut translocation risk | 0
    ICU precautions | 0
    patient monitoring | 0
    infection control measures | -192
    antifungal combination use | 