28 years old | 0
African-woman | 0
gravida 3 | 0
para 0 | 0
past medical history of one miscarriage | -672
past medical history of two abortions | -672
asymptomatic uterine leiomyomas | -672
spontaneous abortion | -336
fever | -336
pelvic pain | -336
vital signs showed a temperature of 38°C | 0
pulse rate of 105/min | 0
blood pressure of 13.3/9.3 kPa | 0
respiratory rate of 16/min | 0
offensive vaginal loss | 0
abdominal tenderness | 0
painful palpation of a large myoma | 0
raised C-reactive protein of 368 mg/L | 0
raised white cell count at 17 × 10^9/L | 0
anemia with Haemoglobin of 95 g/L | 0
platelets at 549 × 10^9/L | 0
PT time at 68% | 0
blood cultures were negative | 0
ultrasonography demonstrated a significant heterogenous leiomyoma | 0
endometrial thickness of 10 mm | 0
contrast enhanced computed tomography (CT) scan | 0
large pelvic mass measuring 16 × 18 × 17 cm | 0
air and heterogeneous tissue suggesting necrosis of a uterine fibroid | 0
three additional masses in the right lumbar region and iliac fossa | 0
free intraperitoneal fluid in the right lumbar region and right iliac fossa | 0
provisional diagnosis of endometritis | 0
conservative treatment with broad spectrum antibiotics | 0
Amoxicillin/clavulanic acid 1 g three times per day | 0
Ofloxacin 400 mg two times per day | 0
deterioration of the patient’s clinical status | 240
persistent fever | 240
persistence of biological inflammatory syndrome | 240
occurrence of bleeding disorders | 240
cholestasis | 240
electrolyte disorders with persistent hypokaliemia | 240
transfer to the intensive care unit | 240
repeat CT scan | 240
persistence of an aspect of reshapes of the necrobiotic myoma complicated with an abscess | 240
exploratory laparotomy | 264
500 mL of a thick reddish-brown fluid | 264
multiple myomas | 264
selective myomectomy of a large myoma of 17 × 15 × 11 cm | 264
padding and hemostatic knots were made using a Vicryl suture | 264
extensive lavage of the peritoneal cavity with warm normal saline | 264
IV antibiotic treatment with Tazocilline, Metronidazole and Amikacin | 264
culture of the peritoneal fluid yielded no growth of bacteria | 264
histopathologic examination of the fibroid revealed a leiomyoma with advanced ischemic necrosis, inflammation and foci of abscess formation | 264
resumption of regular and normal menses | 720
pain had completely resolved | 720
pelvic ultrasound showed an increased volume of the uterus with the largest fibroid measuring 10 cm | 720
spontaneous conception | 17520
fetal growth was normal | 17520
anterior placenta praevia | 17520
cesarean section | 17520
adhesions on the anterior wall of the uterus | 17520
corporeal hysterotomy | 17520
3320 g baby delivered with Apgar’s of 10 | 17520
post-operative recovery was unremarkable | 17520