33 years old | 0
male | 0
admitted to the hospital | 0
general weakness | -744
acute myeloid leukemia | -744
induction chemotherapy | -744
cytarabine | -744
idarubicin | -744
complete remission | -744
consolidation chemotherapy | -744
severe headache | -31
leukemia relapse | -31
intrathecal injection of methotrexate | -31
allogeneic peripheral blood SCT | 0
renal stones | -672
hydronephrosis | -672
busulphan | -4
cyclophosphamide | -4
tacrolimus | -4
methotrexate | -4
micafungin | -4
itraconazole | 0
nonoliguric acute renal failure | 0
discharged | 27
right flank pain | 74
abdominal ultrasonography | 74
non-contrast-enhanced abdominal CT | 74
febrile episode | 75
blood culture | 75
sputum culture | 75
urine culture | 75
PCR for cytomegalovirus | 75
Aspergillus galactomannan antigen | 75
cefepime | 75
amphotericin B deoxycholate | 75
fever subsided | 77
ESWL | 77
cumulative dose of amphotericin B deoxycholate | 96
headache | 96
right flank pain | 96
magnetic resonance imaging of the brain | 96
leptomeningeal leukemic infiltration | 96
CSF cytology | 96
abdominal CT | 96
ureteroscopic lithotripsy | 96
ureteral stent placement | 96
right flank pain subsided | 96
fever developed | 100
abdominal CT | 100
subcapsular hematoma | 100
abscess-like lesion | 100
emergency radical nephrectomy | 109
ruptured area in the right kidney | 109
fungal hyphae | 109
vascular invasion | 109
renal aspergillosis | 109
meropenem | 109
vancomycin | 109
amphotericin B deoxycholate | 109
voriconazole | 109
sepsis progression | 113
died | 113