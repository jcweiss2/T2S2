5-year-old | 0
Chinese | 0
woman | 0
presented to the emergency department | 0
cough | -336
fever | -120
headache | -24
vomiting | -24
altered interactions with her parents | -24
admitted to the pediatric intensive care unit | 0
uncomplicated birth | -26208
normal growth during the first 3 years | -26208
retarded height growth | -17520
decreased activity | -17520
no history of medication | 0
height 109 cm | 0
weight 22 kg | 0
temperature 38.7°C | 0
heart rate 105 beats per minute | 0
respiratory rate 35 breaths per minute | 0
blood pressure 90/55 mmHg | 0
oxyhemoglobin saturation 90% | 0
generalized puffiness | 0
non-pitting edema | 0
capillary refill time >3 seconds | 0
rales | 0
normal cardiac auscultation | 0
soft abdomen | 0
mildly distended abdomen | 0
normal bowel sounds | 0
slightly confused | 0
could not properly respond to commands | 0
hemoglobin 97 g/L | 0
white blood cell count 2.5×10⁹/L | 0
neutrophils 70% | 0
blood platelet 75×10⁹/L | 0
normal electrolytes | 0
normal glucose | 0
normal albumin | 0
normal creatine kinase | 0
normal blood gas | 0
chest CT scan | 0
left lobe pneumonia | 0
mild pleural effusion | 0
echocardiogram | 0
mild pericardial effusion | 0
normal cardiac ejection fraction | 0
MRI scan of the brain | 0
normal cerebrospinal fluid exam | 0
pneumonia | 0
sepsis | 0
empiric antibiotic therapy | 0
immunoglobulin supply | 0
IVIG 2 g/kg | 0
restricted fluid administration | 0
mental status deteriorated | 24
became comatose | 24
temperature dropped to 35°C | 24
developed hypotension | 24
developed arrhythmia | 24
hypoxia | 24
SaO2 decreased to 75% | 24
prolonged Q–T interval | 24
thyroid studies ordered | 0
T4 undetectable | 24
TSH >150 uIU/mL | 24
elevated anti-TPO-Ab | 48
elevated anti-TgAb | 48
thyroid ultrasound | 48
mild bilateral enlargement | 48
small tubercles in the left side | 48
diagnosed with myxedema coma | 24
untreated hypothyroidism | 24
autoimmune thyroiditis | 24
Hashimoto's thyroiditis | 24
intravenous dexamethasone | 24
oral levothyroxine | 24
nasogastric tube | 24
vasopressor | 24
mechanical ventilation | 24
continuous renal replacement treatment | 24
hypotension | 24
hypoxemia | 24
anuria | 24
consciousness restored | 48
temperature returned to normal | 48
extubated | 120
dosage of levothyroxine reduced | 336
discharged | 336
height increased 9 cm | 5832
more active | 5832
father with Hashimoto's thyroiditis | 0
grandmother with Hashimoto's thyroiditis | 0
