61 years old|0
male|0
admitted to the emergency department|0
COVID-19 pneumonia diagnosis|-2160
persistent cough|-2160
expectoration|-2160
streaky hemoptysis|-168
massive hemoptysis|0
respiratory distress|0
low oxygen saturation|0
prior admission for severe COVID-19 pneumonia|-2160
received intravenous methylprednisolone|-2160
received remdesivir|-2160
received tocilizumab|-2160
received prophylactic subcutaneous enoxaparin|-2160
received high flow nasal oxygen|-2160
elevated CRP|-2160
elevated D-dimer|-2160
diabetic|0
bilateral fibrotic sequelae of COVID pneumonia|0
cavitary areas in right lung|0
tested negative for COVID-19 pneumonia|0
shifted to Respiratory intensive treatment unit|0
administered tranexamic acid|0
put on Bilevel Positive Airway Pressure|0
transfused with packed red blood cells|0
CT Pulmonary Angiogram|0
pulmonary arterial pseudoaneurysm|0
alveolar hemorrhage|0
fibro-reticular changes|0
emergency endovascular embolization|0
femoral vein access|0
pulmonary angiogram|0
contrast spill into tracheo-bronchial tree|0
embolisation with coils|0
no further hemoptysis|336
improved oxygen saturation|336
ruled out fungal infection|336
ruled out tuberculosis|336
follow-up CT confirmed successful embolization|336
