66 years old | 0
female | 0
prior TIA | -87600
urea cycle disorder | -87600
elevated amino acids detected on urinalysis | -87600
OTC deficiency confirmed via genetic testing | -87600
admitted in 2016 | -17520
confusion | -17520
gait disturbance | -17520
facial droop | -17520
negative stroke evaluation | -17520
brain MRI no acute changes | -17520
brain toxicity secondary to increased ammonia level | -17520
encephalopathy | -17520
hepatic encephalopathy (HE) signs: inversion of sleep pattern | -17520
mild confusion | -17520
lethargy | -17520
personality changes | -17520
asterixis | -17520
hallucinations | 0
worsening ataxia | 0
fall | 0
abdominal pain | 0
lower-extremity lymphedema | 0
elevated ammonia level of 97 mcg/dL | 0
hypoglycemia | 0
hemoglobin drop from 10 to 8 g/dL | 0
admission | 0
hypotension | 0
seizures | 0
Lorazepam 0.5 mg dose | 0
blood pressure 99/45 mmHg | 0
normal saline bolus | 0
transfer to ICU | 0
blood pressure improved with 500 cc albumin | 0
responsive | 0
Raviciti 1.1 g/mL | 0
lactulose | 0
hyperammonemia | 0
vasopressors | 0
nosocomial pneumonia | 0
secondary septic shock | 0
worsening respiratory status | 0
intubation | 0
vasopressor support | 0
fluctuating ammonia levels between 50 and 170 mcg/dL | 0
fluctuating mental status | 0
glucose levels 40 to 54 mg/dL | 0
D5 infusion | 0
D10 infusion | 0
D20 infusion | 0
normal saline infusion | 0
HAHI syndrome suspected | 0
genetic testing for GLUD-1 gene mutation | 0
elevated alpha-keto glutarate | 0
asymptomatic from elevated ammonia by-products | 0
persistent hypoglycemia | 0
mentation improvement with balanced treatment | 0
dextrose 20 infusion 500 mL/hr | 0
low-protein restricted diet | 0
Raviciti continuation | 0
attempts to wean off dextrose solution | 0
GLUD-1 gene mutation confirmed | 0
decreased GDH levels | 0
elevated alpha-ketoglutarate on urinalysis | 0
Diazoxide use | 0
recurrent hypoglycemia prevention | 0
hyperammonemia prevention |6
adequate nutrition | 0
discharged | 0
