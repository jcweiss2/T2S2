50 years old | 0
female | 0
admitted to the hospital | 0
chronic myeloid leukemia | -1848
blast-phase chronic myeloid leukemia | -528
diagnosed with CML | -1848
treatment with imatinib | -1848
imatinib for 3 months | -1848
progressive disease | -1200
myeloid blastic transformation | -1200
7+3 induction chemotherapy | -1200
intubated | -1200
severe pneumonia | -1200
sepsis | -1200
ICU stay for ~2 months | -1200
bone marrow biopsy | -1200
complete remission | -1200
referred for allo-SCT | -1200
febrile | 0
peripheral blood cultures | 0
central venous port blood cultures | 0
KP susceptible only to tigecycline | 0
venous port infection suspected | 0
venous port removed | 0
treated with tigecycline | 0
treated with meropenem | 0
treatment discontinued after 14 days | 336
in good condition | 336
preparations for allo-SCT | 336
new onset fever | 408
blood cultures revealed KP | 408
same resistance pattern | 408
treated with tigecycline | 408
treated with imipenem | 408
fever resolved | 408
acute-phase parameters returned to normal | 408
treatment discontinued after 2 weeks | 480
fever shortly after | 480
repeated blood cultures | 480
pan-resistant KP | 480
rectal swabs negative for CRKP carrier state | 0
transthoracic echocardiogram | 480
enlarged right cardiac chambers | 480
moderate tricuspid valve insufficiency | 480
mass on tricuspid valve | 480
septic vegetation | 480
tricuspid valve endocarditis diagnosis | 480
operated for excision of vegetation | 480
tricuspid valve repair | 480
treated with imipenem-cilastatin | 480
treated with gentamicin | 480
treated with sulbactam | 480
treatment for 4 weeks | 480
treated for CML with nilotinib | 480
PCR for Bcr/Abl positive | 480
residual disease | 480
infection resolved | 480
allo-SCT performed | 480
neutrophil engraftment on day +15 | 480
thrombocyte engraftment on day +14 | 480
complete remission | 480
complete chimerism | 480
no GVHD | 480
PCR of Bcr/Abl negative | 480
no residual disease | 480
