2-year-old | 0  
    boy | 0  
    father had fever | -672  
    father had exanthema | -672  
    contact with two dogs | -672  
    first symptom was sudden fever (38 °C/١٠٠.٤ °F) | -936  
    received nimesulide | -936  
    received amoxicilin | -936  
    pallor | -912  
    blood test performed | -912  
    leucopenia (2,100 cel/μL) | -912  
    anemia (hemoglobin 8.9 g/dL) | -912  
    thrombocytopenia (75 x103/mL) | -912  
    admitted to the hospital | -888  
    hypoalbuminemia (2.9 g/dL) | -864  
    high AST (1333 U/L) | -864  
    high ALT (972 U/L) | -864  
    high alkaline phosphatase (753 U/L) | -864  
    high LDH (1,714 U/L) | -864  
    prolonged PT (16.6 s) | -864  
    prolonged PTT (54.5 s) | -864  
    hyponatremia (126 mEq/L) | -864  
    elevated C reactive protein (2.4 mg/dL) | -864  
    multiple enlarged lymph nodes in the neck | -864  
    hepatomegaly (4 cm) | -864  
    splenomegaly (5 cm) | -864  
    erythematous macular non%itching rash on thorax thighs and buttocks | -864  
    single left inguinal adenopathy | -864  
    fever with nocturnal and needle pattern | -864  
    coughs without consolidations or pneumonia | -864  
    bone marrow aspiration performed | -864  
    activated lymphocytes without leukemia | -864  
    persistence of cytopenia | -864  
    anemia (Hb 6.3 g/dL) | -864  
    deep neutropenia (0.3 x103/μL) | -864  
    thrombocytopenia (98x103/mL) | -864  
    normal kidney function | -864  
    hemorrhagic syndrome | -864  
    managed with transfusions | -864  
    persistent hyponatremia (126-128 mEq/L) | -864  
    liver failure with incoagulable PT | -864  
    persistent hypoalbuminemia | -864  
    LDH peaked over 6700 UI/L | -864  
    serological tests performed (HIV, Epstein-Barr, Hepatitis A, B, C, Toxoplasma, cytomegalovirus, rubella, herpes, Treponema) | -864  
    Weil-Felix reactions | -864  
    all tests negative | -864  
    bone marrow biopsy with cellularity 70% | -672  
    myeloid-erythroid ratio inverted | -672  
    myeloid hypoplasia | -672  
    erythroid series hyperplasia with megaloblastic maturation | -672  
    megakaryocytic series hypolobulated nuclei | -672  
    histiocytes with hemophagocytosis | -672  
    䋼 lymph node biopsy with histiocytic infiltration | -672  
    immunohistochemistry for Langerhans ruled out | -672  
    radiographs ruled out Langerhans disease | -672  
    jaundice developed | -504  
    doxycycline initiated (2.2 mg/kg/day) | -504  
    fever remission within 48 hours | -480  
    improvement of general condition | -480  
    new fever peaks | -480  
    jaundice reappeared | -480  
    asthenia reappeared | -480  
    increased triglycerides | -480  
    persistence of cytopenia | -480  
    low fibrinogen levels | -480  
    Leptospira interrogans ruled out by PCR | -480  
    splenomegaly confirmed | -480  
    diagnosis of HLH | -480  
    started methylprednisolone (30 mg/kg/day) | -480  
    nested PCR for Rickettsia 17-kDA gene negative | -480  
    indirect immunofluorescence assay for IgM and IgG (Rickettsia rickettsii and R. typhi) | -480  
    negative result on day 14 | -480  
    seroconversion on day 27 (IgM 1:128, IgG 1:512 to R. typhi) | -480  
    hemorrhagic syndrome with petechiae and gingivorrhagia | -336  
    admitted to Pediatric ICU | -336  
    neurological deterioration | -336  
    respiratory deterioration | -336  
    meropenem | -336  
    vancomycin | -336  
    amphotericin B | -336  
    nosocomial sepsis suspected | -336  
    blood cultures negative | -336  
    doxycycline suspended | -336  
    gastric bleeding | -336  
    dexamethasone added | -336  
    poor response | -336  
    abdominal ultrasound with hepatic and kidney damage | -336  
    ascites reported | -336  
    urine output decreased | -336  
    neurological worsening | -336  
    hemodynamic worsening | -336  
    mechanical ventilation started | -336  
    vasopressors started | -336  
    alveolar diffuse hemorrhage | -336  
    anuria developed | -336  
    died | 0  
    post-mortem lymph node biopsy | 24  
    IHC positive for Rickettsia | 24  
    <|eot_id|>
    2-year-old | 0  
    boy | 0  
    father had fever | -672  
    father had exanthema | -672  
    contact with two dogs | -672  
    first symptom was sudden fever (38 °C/١٠٠.٤ °F) | -936  
    received nimesulide | -936  
    received amoxicilin | -936  
    pallor | -912  
    blood test performed | -912  
    leucopenia (2,100 cel/μL) | -912  
    anemia (hemoglobin 8.9 g/dL) | -912  
    thrombocytopenia (75 x103/mL) | -912  
    admitted to the hospital | -888  
    hypoalbuminemia (2.9 g/dL) | -864  
    high AST (1333 U/L) | -864  
    high ALT (972 U/L) | -864  
    high alkaline phosphatase (753 U/L) | -864  
    high LDH (1,714 U/L) | -864  
    prolonged PT (16.6 s) | -864  
    prolonged PTT (54.5 s) | -864  
    hyponatremia (126 mEq/L) | -864  
    elevated C reactive protein (2.4 mg/dL) | -864  
    multiple enlarged lymph nodes in the neck | -864  
    hepatomegaly (4 cm) | -864  
    splenomegaly (5 cm) | -864  
    erythematous macular non%itching rash on thorax thighs and buttocks | -864  
    single left inguinal adenopathy | -864  
    fever with nocturnal and needle pattern | -864  
    coughs without consolidations or pneumonia | -864  
    bone marrow aspiration performed | -864  
    activated lymphocytes without leukemia | -864  
    persistence of cytopenia | -864  
    anemia (Hb 6.3 g/dL) | -864  
    deep neutropenia (0.3 x103/μL) | -864  
    thrombocytopenia (98x103/mL) | -864  
    normal kidney function | -864  
    hemorrhagic syndrome | -864  
    managed with transfusions | -864  
    persistent hyponatremia (126-128 mEq/L) | -864  
    liver failure with incoagulable PT | -864  
    persistent hypoalbuminemia | -864  
    LDH peaked over 6700 UI/L | -864  
    serological tests performed (HIV, Epstein-Barr, Hepatitis A, B, C, Toxoplasma, cytomegalovirus, rubella, herpes, Treponema) | -864  
    Weil-Felix reactions | -864  
    all tests negative | -864  
    bone marrow biopsy with cellularity 70% | -672  
    myeloid-erythroid ratio inverted | -672  
    myeloid hypoplasia | -672  
    erythroid series hyperplasia with megaloblastic maturation | -672  
    megakaryocytic series hypolobulated nuclei | -672  
    histiocytes with hemophagocytosis | -672  
    lymph node biopsy with histiocytic infiltration | -672  
    immunohistochemistry for Langerhans ruled out | -672  
    radiographs ruled out Langerhans disease | -672  
    jaundice developed | -504  
    doxycycline initiated (2.2 mg/kg/day) | -504  
    fever remission within 48 hours | -480  
    improvement of general condition | -480  
    new fever peaks | -480  
    jaundice reappeared | -480  
    asthenia reappeared | -480  
    increased triglycerides | -480  
    persistence of cytopenia | -480  
    low fibrinogen levels | -480  
    Leptospira interrogans ruled out by PCR | -480  
    splenomegaly confirmed | -480  
    diagnosis of HLH | -480  
    started methylprednisolone (30 mg/kg/day) | -480  
    nested PCR for Rickettsia 17-kDA gene negative | -480  
    indirect immunofluorescence assay for IgM and IgG (Rickettsia rickettsii and R. typhi) | -480  
    negative result on day 14 | -480  
    seroconversion on day 27 (IgM 1:128, IgG 1:512 to R. typhi) | -480  
    hemorrhagic syndrome with petechiae and gingivorrhagia | -336  
    admitted to Pediatric ICU | -336  
    neurological deterioration | -336  
    respiratory deterioration | -336  
    meropenem | -336  
    vancomycin | -336  
    amphotericin B | -336  
    nosocomial sepsis suspected | -336  
    blood cultures negative | -336  
    doxycycline suspended | -336  
    gastric bleeding | -336  
    dexamethasone added | -336  
    poor response | -336  
    abdominal ultrasound with hepatic and kidney damage | -336  
    ascites reported | -336  
    urine output decreased | -336  
    neurological worsening | -336  
    hemodynamic worsening | -336  
    mechanical ventilation started | -336  
    vasopressors started | -336  
    alveolar diffuse hemorrhage | -336  
    anuria developed | -336  
    died | 0  
    post-mortem lymph node biopsy | 24  
    IHC positive for Rickettsia | 24  
    
