33 years old | 0
male | 0
admitted to the intensive care unit | 0
severe hypotension | 0
persistent fever | 0
dyspnea | 0
chest pain | 0
diarrhea | 0
blood pressure of 47/29 mmHg | 0
tachycardia | 0
need for oxygen therapy | 0
hepatojugular reflux | 0
cardiogenic shock | 0
bilateral conjunctivitis | 0
cheilitis | 0
hypertension | -4032
fever episode lasting for 5 days | -4032
myalgia | -4032
dysgeusia | -4032
anosmia | -4032
COVID-19 | -4032
leukocytosis | 0
normocytic anemia | 0
elevated liver enzyme levels | 0
elevated creatine kinase levels | 0
acute kidney injury | 0
elevated CRP levels | 0
elevated brain natriuretic peptide levels | 0
elevated D-dimer levels | 0
elevated troponin levels | 0
sinus tachycardia | 0
TTE showing global hypokinesis | 0
dilated inferior vena cava | 0
reduced ejection fraction | 0
acute myocarditis | 0
high titers of SARS-CoV-2 IgG | 0
multiple coronary aneurysms | 336
hemodynamic support | 0
norepinephrine infusion | 0
dobutamine infusion | 0
IVIG | 0
prednisone | 0
aspirin | 0
resolution of symptoms by day 10 | 240
CRP levels dropped to 10 mg/l | 240
control TTE showing normal left ventricular function | 168
cardiac magnetic resonance imaging unremarkable | 168
discharged | 288
partial regression of coronary aneurysms | 1344
normalization of left ventricular function | 1344
complete disappearance of all aneurysms | 3600
