83 years old | 0
female | 0
insulin-dependent diabetes mellitus | 0
hypertension | 0
hyperlipidemia | 0
diastolic heart failure | 0
diabetic gastroparesis | 0
chronic kidney disease | 0
nausea | -72
substernal epigastric abdominal discomfort | -72
belching | -72
poor oral intake | -72
mild right upper quadrant tenderness | 0
aperistalsis of the esophageal body | 0
elevated LES pressure | 0
type I achalasia | 0
decreased motility of the esophagus | 0
BT injections | 0
immediate improvement in symptoms | 0
right shoulder pain | 504
NSAIDS for pain relief | 504
intra-articular steroid injections | 504
persistent symptoms | 504
white blood cell count of 30.7 K/μL | 522
CT scan of the abdomen | 522
5.8 cm x 6.9 cm x 2.3 cm fluid collection | 522
vancomycin and piperacillin/tazobactam | 522
abscess drainage | 522
fluid cultures grew Streptococcus intermedius | 522
vancomycin trough after the third dose was 32 μg/ml | 522
discontinuation of vancomycin and piperacillin/tazobactam | 522
ampicillin/sulbactam 3 g every 12 hours | 522
leukocytosis improvement | 522
interval decrease in abscess size | 522
generalized edema | 522
acute kidney injury | 522
hemodialysis initiation | 522
unresponsive | 528
endotracheal intubation | 528
septic shock | 528
vasopressor support | 528
antibiotics escalation to meropenem and vancomycin | 528
ischemic hepatopathy | 528
large left pleural effusion | 528
chest tube placement | 528
atrial fibrillation with rapid ventricular response | 528
comfort care measures | 480
death | 504