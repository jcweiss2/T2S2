57 years old | 0
male | 0
lepromatous leprosy | -720
treatment with rifampicin/clofazimine/dapsone | -720
abdominal distension | 0
constipation | 0
vomiting | 0
10-kg weight loss | 0
peripheral lymphadenopathy | 0
distended abdomen | 0
positive shifting dullness | 0
mural thickening of the terminal ileum | 0
enlarged mesenteric lymph nodes | 0
mesenteric fat stranding | 0
intra-abdominal free fluid | 0
abdominal granulomatous infection | 0
neoplastic process | 0
abdominal paracentesis | 0
atypically large lymphocytes | 0
high-grade lymphoma | 0
flow cytometry | 0
abnormal CD4/CD8 double-negative T-cell population | 0
cervical lymph node biopsy | 0
high-grade peripheral T-cell lymphoma | 0
bone marrow examination | 0
no involvement of T-cell NHL | 0
stage IV lymphoma | 0
dexamethasone | 0
tumor-lysis syndrome precautions | 0
severe sepsis | 24
transfer to ICU | 24
antibiotics | 24
antifungals | 24
ICU care | 24
recovered | 168
transfer to national cancer center | 168
EPOCH chemotherapy protocol | 168
CNS prophylaxis | 168
intrathecal methotrexate | 168
febrile neutropenia episodes | 336
recurrent bacteremia | 336
generalized weakness | 336
no sensory changes | 336
no clear fatigability | 336
decreased power in proximal and distal muscles | 336
normal distal latencies | 336
normal compound muscle action potential | 336
normal conduction velocities | 336
normal F waves | 336
normal sensory nerve studies | 336
needle electromyogram | 336
poor recruitment effects | 336
repetitive nerve stimulation | 336
significant incremental response | 336
presynaptic neuromuscular junction disorder | 336
LEMS | 336
intravenous immunoglobulins | 336
significant improvement of motor function | 360
ambulate | 360
consolidation by autologous bone marrow transplant | 720
recurrent bacteremia and sepsis | 720
multiorgan failure | 720
death | 1440