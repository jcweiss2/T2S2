65 years old|0
male|0
admitted to the emergency department|0
persistent high-grade fever|-240
nausea|-240
vomiting|-240
generalized weakness|-240
hypertension| -4320
benign prostate hyperplasia| -17520
regular medication for hypertension| -4320
regular medication for benign prostate hyperplasia| -17520
intermittent high-grade fever| -720
vomiting| -720
loss of weight| -720
night-sweats| -720
conscious|0
well-built|0
oriented|0
lethargic|0
febrile temperature of 101 °F|0
mild hepatosplenomegaly|0
conjunctival pallor|0
hepatosplenomegaly|0
fatty liver|0
mild urinary bladder wall thickening|0
mild cystitis|0
mean corpuscular volume: 78 fL|24
absolute neutrophil count: 2.17 × 103/μL|24
microcytic hypochromic anemia|24
hemoglobin: 9.4 g/dL|24
leukocytopenia|24
leukocyte count: 2.94 × 103/μL|24
total platelet count: 90 × 103/μL|24
bicytopenia|24
raised liver transaminases|24
total bilirubin: 0.85 mg/dL|24
serum triglyceride within normal limits|24
plasma fibrinogen levels within normal limits|24
hepatitis B negative|24
hepatitis C negative|24
HIV negative|24
malaria negative|24
dengue negative|24
scrub typhus negative|24
urine culture negative|24
sputum culture negative|24
blood culture negative|24
continuous fever|192
increasing cytopenias|192
fatigue|192
organomegaly|192
bone marrow biopsy|192
trephine biopsy|192
erythroid hyperplasia|192
megaloblastic erythropoiesis|192
erythroid phagocytosis|192
lymphophagocytosis|192
raised lactate dehydrogenase: 1552.30 IU/L|192
hyperferritinemia: >1700 ng/mL|192
hyponatremia: 117 mmol/L|192
decreased total protein: 4.72 g/dL|192
Acid-Fast Bacilli negative|192
MTB detected|192
Rifampicin indeterminate|192
mild hepatomegaly|192
prostatomegaly|192
hepatomegaly|192
external iliac lymphadenopathy|192
disseminated tuberculosis|192
fulfillment of 5 out of 8 HLH diagnostic criteria|360
supportive measures initiated|360
broad-spectrum intravenous antibiotics initiated|360
transfused with two units of PRBC|360
modified Anti-Tubercular Treatment initiated|360
ethambutol|360
levofloxacin|360
streptomycin|360
methylprednisolone|360
Intravenous Immunoglobulin|360
sudden onset breathlessness|384
SpO2 -90%|384
shifted to intensive care unit|384
hemoglobin: 7.7 g/dL|384
leukocyte count: 0.90 × 103/μL|384
total platelet count: 32 × 103/μL|384
Urea: 91 mg/dL|384
LDH: 8000 U/L|384
AST: 1000 U/L|384
creatinine: 1.39 mg/dL|384
ALT: 230 U/L|384
status epilepticus|384
poor Glasgow Coma Scale|384
intubated|384
failed resuscitation|384
death|480
