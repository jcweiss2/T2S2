69 years old | 0
man | 0
coronary artery disease | 0
aspirin | 0
hypertension | 0
type 2 diabetes mellitus | 0
fever | -168
malaise | -168
progressive shortness of breath | -168
temperature of 103.1 °F | 0
pulse of 106 beats per minute | 0
respiratory rate of 18 per minute | 0
blood pressure of 142/70 mm Hg | 0
saturation of 89% on room air | 0
decreased breath sounds bilaterally at base | 0
crepitations | 0
hemoglobin 12.7 g/dL | 0
white blood cell count of 4.5 × 10³ | 0
platelet count of 164 × 10³ | 0
neutrophil 76.4% | 0
lymphocyte 14.9% | 0
absolute lymphocytes 0.7 | 0
C-reactive protein 12.07 mg/dL | 0
D-dimer 570 ng/mL | 0
influenza A and B serology negative | 0
COVID-19 RT-PCR positive | 0
chest X-ray bilateral infiltrates at lung bases | 0
hydroxychloroquine | 0
azithromycin | 0
supplemental oxygen with nasal cannula | 0
enoxaparin 40 mg subcutaneous prophylactic | 0
respiratory condition worsened | 24
repeat chest X-ray worsening bilateral infiltrates | 24
transitioned to optiflow | 24
D-dimer up trended to 1,763 ng/mL | 24
continued on aspirin | 24
therapeutic enoxaparin | 24
abdominal pain | 480
pulse of 113 beats per minute | 480
blood pressure 74/45 mm Hg | 480
hemoglobin level of 8.9 g/dL | 480
hypovolemic shock | 480
CT scan of abdomen and pelvis without contrast | 480
hemorrhage along entire length of right psoas muscle | 480
transferred to ICU | 480
resuscitated with 2 L intravenous fluid | 480
3 units of PRBC | 480
vasopressors | 480
did not respond to fluids | 480
vasopressor requirement increased | 480
post-transfusion hemoglobin of 6.6 g/dL | 480
two more units of PRBC | 480
1 unit of fresh frozen plasma | 480
arterial embolization planned | 480
left common femoral artery accessed | 480
abdominal aortogram performed | 480
subtle extravasation from right L3 and L4 lumbar arteries | 480
selectively catheterized with 5 French Mickelson catheter | 480
high flow microcatheter placed | 480
active extravasation identified | 480
Embosphere particles administered | 480
four 4 mm microcoils | 480
no active contrast extravasation | 480
one more unit of PRBC | 480
hemoglobin stabilized to 7.9 g/dL | 480
vasopressor requirement decreased | 480
vasopressors discontinued | 480
repeat CT scan decreased size of hematoma | 504
remained in ICU | 504
stable hemoglobin level | 504
no further bleeding | 504
weaned off optiflow | 504
transferred to medical floors | 504
