56 years old| 0
male| 0
chronic hepatitis B| -17520
hepatocellular carcinoma| -17520
abdominal distension| -17520
dynamic CT scan of the liver| -17520
five hypervascular lesions| -17520
cirrhosis| -17520
splenomegaly| -17520
esophageal varices| -17520
no ascites| -17520
local treatment with RFA| 0
small ventricular septal defect| 0
left to right shunting| 0
normal chamber sizes| 0
normal left ventricular ejection fraction| 0
Child Class A compensated liver disease| 0
serum albumin 32 g/L| 0
serum bilirubin 21 µmol/L| 0
ALT 45 IU/L| 0
AST 54 IU/L| 0
platelet count 61 × 10^9/L| 0
INR 1.2| 0
AFP 23.8 ng/mL| 0
general anesthesia| 0
fluoroscopic CT guidance| 0
RFA needle placement| 0
tumour ablation| 0
coagulation necrosis| 0
expanding pericardial effusion| 0
hemorrhagic cardiac tamponade| 0
pericardiocentesis| 0
aspiration of 300 mL blood| 0
persistent hypotension| 0
emergency sternostomy| 0
two liters of blood evacuated| 0
puncture wound at anterior cardiac vein| 0
inflammatory changes in adjacent diaphragm|?
repair of anterior cardiac vein| 0
hemostasis secured| 0
post-surgery stability| 24
liver failure| 456
upper gastrointestinal bleeding| 456
pneumonia| 456
sepsis| 456
expiration| 456
no pericardial fluid| 0
no liver abscess| 0
no intraperitoneal hemorrhage| 0
no biloma| 0
no ground pad burn| 0
no diaphragmatic injury| 0
no pneumothorax| 0
no pleural effusion| 0
no bowel perforation| 0
no hepatic infarction| 0
no renal infarction| 0
no tumor seeding| 0
