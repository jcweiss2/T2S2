54 years old | 0
male | 0
admitted to the hospital | 0
weight 168 kg | 0
height 1.75 m | 0
body mass index 56 kg/m2 | 0
chronic obstructive pulmonary disease | -8760
obstructive sleep apnea | -8760
continuous positive airway pressure | -8760
acute renal failure | 0
sepsis | 0
Fournier’s gangrene | 0
emergent debridement | 0
respiratory failure | 0
intubation | 0
metabolic acidosis | 0
coronary artery disease | -8760
percutaneous coronary intervention | -8760
stenting | -8760
30 pack-year smoking history | -8760
morbid obesity | -8760
respiratory distress | 0
tachypnea | 0
diffuse bilateral wheezing | 0
mouth opening of three finger-breadths | 0
Mallampati airway classification 3 | 0
thyromental distance of 6 cm | 0
neck circumference of 44 cm | 0
blood oxygen saturation 99% | 0
fraction of inspired oxygen of 0.5 | 0
cyanotic | 0
blood oxygen saturation ~85% | 0
coarse, low-pitched wheezing | 0
dyspnea | 0
bronchodilators | 0
elevated prothrombin time | 0
international normalized ratio 3.6 | 0
septic shock | 0
regional anesthesia contraindicated | 0
general anesthetic | 0
awake fiberoptic endotracheal intubation | 0
bilateral superior laryngeal nerve block | 0
transtracheal instillation of 4% lidocaine | 0
fiberoptic intubation | 0
tracheomalacia | 0
endotracheal tube insertion | 0
debridement of Fournier’s gangrene | 0
vasoactive agents | 0
phenylephrine | 0
intraoperative arterial blood gas | 0
pH 7.26 | 0
partial pressure of carbon dioxide 34 mmHg | 0
partial pressure of oxygen 320 mmHg | 0
HCO3− levels 16.0 | 0
base excess −11 | 0
blood oxygen saturation 100% | 0
intensive care unit | 0
antibiotics | 0
inotropic support | 0
pressure-regulated volume control ventilation | 0
fraction of inspired oxygen of 1.0 | 0
respiratory rate of 20 breaths per minute | 0
peak inspiratory pressure of 25 mmHg | 0
positive end-expiratory pressure of 7 mmHg | 0
acute respiratory distress syndrome | 24
computed tomography scan of the chest | 24
bilateral infiltrates in lung bases | 24
multiorgan dysfunction | 120
hepatic dysfunction | 120
renal dysfunction | 120
cardiac dysfunction | 120
pulmonary dysfunction | 120
death | 120