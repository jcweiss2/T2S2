62 years old | 0
male | 0
transferred to the emergency department | 0
high fever | 0
39.0°C | 0
dark urine | 0
worsened condition | -2160
repeated dehiscence | -2160
exudation of wounds | -2160
sacrococcygeal region wounds | -2160
lumbar vertebral injury | -262080
paralysis | -262080
sacrococcygeal bedsores | -87600
debridement | -87600
muscle flap application | -87600
infected wound | 0
size 2 × 4 cm | 0
depth reaching sacrum surface | 0
amyotrophy of both lower limbs | 0
disappearance of cutaneous sensation | 0
absence of physiological reaction | 0
absence of pathological character |1 0
CK level significantly elevated | 0
multidisciplinary team consultation | 0
debridement | 24
intraoperative exploration | 24
distal wound debrided | 24
distal wound sutured | 24
pus removed | 24
necrotic muscle removed | 24
fresh granulation tissue observed | 24
frequent dressing changes | 24
antimicrobial therapy | 24
correction of electrolyte imbalances | 24
correction of acidosis | 24
nutritional support | 24
suture area dry | 72
suture area clean | 72
no swelling | 72
no exudation | 72
dark urine lightened | 24
urine normal color | 120
fever resolved | 72
CK peaked | 24
CK decreased | 24
CK returned to normal | 216
white blood cell count decreased | 24
white blood cell count returned to normal | 168
C-reactive protein decreased | 24
C-reactive protein returned to normal | 264
discharged | 720
wound healed | 2160
no sign of infection | 2160
pressure ulcers | 0
rhabdomyolysis | 0
myoglobinuria | 0
acute infection | 0
severe renal dysfunction | 0
metabolic disturbance | 0
multidisciplinary diagnosis and treatment model | 0
anesthesia | 0
thorough debridement | 0
chronic sacrococcygeal pressure ulcers | 0
infection | 0
paraplegia | 0
loss of skin sensation | 0
acute kidney injury risk | 0
sepsis risk | 0
