41 years old | 0
    morbidly obese | 0
    admitted to the hospital | 0
    painful bilateral oedema of lower legs | -24
    generalized abdominal pain | -24
    liver cirrhosis | -24
    excessive alcohol abuse | -24
    hepatitis C infection | -24
    portal hypertension | -24
    oesophageal varices | -24
    febrile (37.6 °C) | 0
    bilateral pitting oedema | 0
    superficial pre-tibial abrasions over left leg | 0
    normal capillary refill time | 0
    distal pulses present in lower limbs | 0
    unremarkable abdominal examination | 0
    unremarkable respiratory examination | 0
    unremarkable cardiovascular examination | 0
    unremarkable neurological examination | 0
    low haemoglobin (11.2 g/dl) | 0
    low platelet count (44 × 10^9/l) | 0
    low albumin (19 g/l) | 0
    elevated bilirubin (36 μmol/l) | 0
    elevated CRP (37 mg/l) | 0
    elevated INR (2.1) | 0
    elevated lactate (8.6 mmol/l) | 0
    liver enzymes at upper limits of normal | 0
    Child's B cirrhosis classification | 0
    blood cultures | 0
    swab of left leg | 0
    intravenous flucloxacillin | 0
    intravenous benzylpenicillin | 0
    suspected cellulitis | 0
    left leg swelling increased | 24
    erythematous skin | 24
    tender skin | 24
    induration | 24
    blistering | 24
    CRP increased (101.7 mg/l) | 24
    intravenous ciprofloxacin | 24
    intravenous cephazolin | 24
    left leg duplex ultrasound | 24
    severe oedema below knee | 24
    knee joint effusion | 24
    no deep vein thrombosis | 24
    CT scan of legs | 24
    bilateral knee joint effusions | 24
    non-specific synovitis | 24
    no necrotizing fasciitis | 24
    blood cultures grew A. baumannii | 48
    multi-drug resistance to amoxicillin | 48
    multi-drug resistance to amoxicillin/clavulanate | 48
    multi-drug resistance to ceftriaxone | 48
    multi-drug resistance to ceftazidime | 48
    sensitivity to co-trimoxazole | 48
    sensitivity to gentamycin | 48
    sensitivity to meropenem | 48
    sensitivity to ciprofloxacin | 48
    sensitivity to ticarcillin/clavulanate | 48
    antibiotic regime changed to meropenem | 48
    antibiotic regime changed to vancomycin | 48
    conservative management with leg elevation | 48
    conservative management with compression bandages | 48
    referred to reconstructive surgeons | 48
    referred to orthopaedic surgeons | 48
    evaluation for septic arthritis | 48
    evaluation for compartment syndrome | 48
    exclusion of necrotizing fasciitis | 48
    MRI scan of lower legs | 72
    extensive subcutaneous oedema left leg | 72
    moderate subcutaneous oedema right leg | 72
    bilateral joint effusions | 72
    cellulitic changes left leg | 72
    extensive myositis left leg | 72
    possible fasciitis | 72
    suspicion of compartment syndrome | 72
    no immediate surgical intervention | 72
    left leg erythematous | 72
    left leg bullous | 72
    left leg blistering | 72
    added lincomycin | 72
    spiked fever (38.4 °C) | 96
    left leg surgically explored | 96
    general anaesthesia | 96
    leg tourniquet applied | 96
    longitudinal incision | 96
    no necrotizing fasciitis found | 96
    no compartment syndrome found | 96
    no abscess | 96
    no drainable collection | 96
    extensive subcutaneous oedema | 96
    circumferential debridement of fat necrosis | 96
    circumferential debridement of muscle | 96
    washout of left leg wound | 96
    VAC dressing applied | 96
    antibiotics continued | 96
    subcutaneous fat sent for culture | 96
    fascia sent for culture | 96
    histopathological review | 96
    cultures confirmed A. baumannii | 96
    remained ventilated post-operatively | 96
    commenced noradrenaline infusion | 96
    hypotension | 96
    cultures resistant to amoxicillin | 96
    cultures resistant to augmentin | 96
    cultures resistant to ceftriaxone | 96
    cultures resistant to ceftazidime | 96
    cultures sensitive to co-trimoxazole | 96
    cultures sensitive to gentamicin | 96
    antibiotic regime changed to ciprofloxacin | 96
    antibiotic regime changed to meropenem | 96
    antibiotic regime changed to lincomycin | 96
    vancomycin ceased | 96
    further surgical debridement | 168
    necrotic circumferential subcutaneous fat | 168
    circumferential debridement performed | 168
    extensive washout with hydrogen peroxide | 168
    new VAC dressing applied | 168
    histopathology revealed epidermal infarction | 168
    histopathology revealed dermal infarction | 168
    focal fat necrosis | 168
    acute inflammation | 168
    no histological evidence of fasciitis | 168
    tailored antibiotics to meropenem | 168
    tailored antibiotics to ciprofloxacin | 168
    two further surgical procedures | 312
    VAC dressing changed | 312
    wound clean | 312
    areas of necrosis along wound edges | 312
    minor debridement | 312
    VAC dressing replaced | 312
    VAC dressing replaced again | 384
    significant wound improvement | 384
    small areas of necrotic tissue | 384
    necrotic tissue attached to fascia | 384
    viable musculature | 384
    minor debridement performed | 384
    removal of necrotic tissue | 384
    removal of fascia | 384
    samples sent for microscopy | 384
    wound washed with hydrogen peroxide | 384
    jaundice | 672
    worsening hepatic function | 672
    worsening renal function | 672
    condition deterioration | 672
    developed hepatic failure | 672
    developed circulatory failure | 672
    developed respiratory failure | 672
    developed haematological failure | 672
    blood glucose fluctuations | 672
    inotrope dependency | 672
    single glucose reading of 10 mmol/l | 672
    insulin required | 672
    required vasopressor support | 504
    significant tissue loss in lower limbs | 504
    decision to palliate | 504
    death | 504