22 years old | 0
    male | 0
    admitted to the hospital | 0
    intermittent fevers | -336
    headache | -336
    fatigue | -336
    malaise | -336
    nausea | -336
    vomiting | -336
    occasional episodes of diarrhea | -336
    nosebleeds | -336
    non-productive cough | -336
    sore throat | -336
    headache associated with light sensitivity | -336
    rash began over thighs | -72
    rash spread to entire body | -72
    no shortness of breath | 0
    no chest pain | 0
    no bloody stools | 0
    no neck stiffness | 0
    working as a taxidermist | -72
    cat at home | 0
    two dogs at home | 0
    possible fleas | 0
    unconfirmed rats in home | 0
    afebrile | 0
    blood pressure 97/47 | 0
    pulse rate 136 bpm | 0
    respiratory rate 22 bpm | 0
    petechial rash on trunk | 0
    petechial rash on upper extremities | 0
    petechial rash on lower extremities | 0
    no nuchal rigidity | 0
    hyponatremia (sodium 126 mmol/L) | 0
    elevated BUN (111 mg/dL) | 0
    elevated creatinine (3.14 mg/dL) | 0
    elevated AST (421 U/L) | 0
    elevated ALT (135 U/L) | 0
    elevated ALP (158 U/L) | 0
    elevated D-dimer (17.55 µg/mL) | 0
    low fibrinogen (94 mg/dL) | 0
    elevated lactic acid (2.34 mmol/L) | 0
    thrombocytopenia (35,000/mm³) | 0
    elevated WBC (13,830/mm³) | 0
    diagnosed with severe sepsis | 0
    diagnosed with DIC | 0
    admitted to MICU | 0
    vancomycin treatment | 0
    ceftriaxone treatment | 0
    lumbar puncture not performed due to thrombocytopenia | 0
    stabilized | 24
    seen by infectious diseases specialist | 24
    differential diagnosis: viral infection | 24
    differential diagnosis: ehrlichiosis | 24
    differential diagnosis: murine typhus | 24
    EBV serology negative | 24
    parvovirus serology negative | 24
    Ehrlichial DNA assay negative | 24
    Rickettsia typhi titers requested | 24
    Rickettsia typhi IgM and IgG positive | 48
    vancomycin changed to doxycycline | 24
    hematology consultation | 24
    cryoprecipitate administration | 24
    no schistocytes on blood smear | 24
    DIC excluded | 24
    fever resolved | 72
    hemodynamically stable for transfer | 72
    repeat infection work-up | 120
    high Rickettsia typhi IgM (1:2048) | 120
    high Rickettsia typhi IgG (1:512) | 120
    oral doxycycline 100 mg twice daily | 120
    discharged after improvement | 168
    
    
    