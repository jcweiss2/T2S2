21 years old | 0
male | 0
Prader-Willi syndrome | -7560
neonatal hypotonia | -7560
distinctive facial features | -7560
poor growth in infancy | -7560
hyperphagia | -6840
severe obesity | -6840
short stature | -6840
hypogonadism | -6840
intellectual disability | -6840
behavior problems | -6840
birth weight 3.3 kg | -7560
gestational age 39 weeks | -7560
cesarean section | -7560
poor feeding | -7560
bilateral undescended testicles | -7560
obesity | -5760
hyperphagia | -5760
diagnosed with PWS | -5760
methylation polymerase chain reaction | -5760
height 151 cm | -5760
weight 75 kg | -5760
recombinant growth hormone treatment | -5760
methylphenidate | -5760
attention deficit hyperactivity disorder | -5760
polysomnography | -5760
obstructive sleep apnea | -5760
tonsillectomy | -5040
gonadotropin-releasing hormone deficiency | -4320
growth hormone deficiency | -4320
uncontrolled glycemic status | -4320
osmotic symptoms | -4320
polyuria | -4320
polydipsia | -4320
polyphagia | -4320
diagnosed with DM | -4320
metformin | -4320
glipizide | -3600
long-acting insulin | -3600
oxygen saturation 50% | -3600
positive pressure ventilation | -3600
poor compliance | -3600
normal ventricle size | -3600
normal systolic function | -3600
dyspnea | 0
loss of consciousness | 0
height 164 cm | 0
weight 185.7 kg | 0
BMI 69.04 kg/m2 | 0
blood pressure 96/25 mmHg | 0
body temperature 39℃ | 0
heart rate 93 beats per minute | 0
respiratory rate 28 per minute | 0
oxygen saturation 63% | 0
periorbicular cyanosis | 0
respiratory distress | 0
skin ulcers | 0
macular rash | 0
cardiomegaly | 0
haziness in the right lung | 0
arterial blood gas analysis | 0
pH 6.9 | 0
PCO2 147 | 0
PO2 72.1 | 0
HCO3 29.3 | 0
intubation | 0
synchronized intermittent mandatory ventilation | 0
hemoglobin level 15 g/dL | 0
white blood cell level 19,620/μL | 0
erythrocyte sedimentation rate 49 mm/hr | 0
C-reactive protein 2.37 mg/dL | 0
lactic acid 10.37 mmol/L | 0
albumin 3.8 g/dL | 0
aspartate aminotransferase/alanine aminotransferase 51 U/L/59 U/L | 0
blood urea nitrogen/creatinine 34.9 mg/dL/0.93 mg/dL | 0
fasting glucose level 141 mg/dL | 0
glycosylated hemoglobin 8.2% | 0
thyroid stimulating hormone/free T4 2.576 uIU/mL/1.01 ng/dL | 0
Troponin I level 0.844 ng/mL | 0
creatine kinase-MB 3.73 ng/mL | 0
pro-B-type natriuretic peptide 1,904 pg/mL | 0
normal saline | 0
noradrenalin | 0
cefotaxime | 0
midazolam | 0
fentanyl | 0
physiotherapy | 0
transesophageal echocardiography | 0
dilated RV cavity | 0
decreased RV systolic function | 0
pulmonary hypertension | 0
right heart failure | 0
cor pulmonale | 0
furosemide | 0
caloric restriction | 0
skin care | 0
rehabilitation | 0
pressure-relieving mattress | 0
weighing machine | 0
clindamycin | 96
wound dressing | 96
total parenteral nutrition | 96
ventilator mode change | 168
pressure-control SIMV | 168
weight loss 5.8 kg | 240
pulmonary congestion | 240
pleural effusion | 240
target balance of I/O -1,500–2,000 mL/day | 240
weight loss 1.8 kg per day | 240
lung congestion improvement | 240
enteral nutrition | 336
nasogastric tube | 336
insulin injections | 336
full enteral feeding | 504
oral feeding | 588
discharge | 588
weight 131.4 kg | 588
BMI | 588
furosemide 0.3 mg/kg/day | 588
spironolactone 0.19 mg/kg/day | 588
metformin 15.2 mg/kg/day | 588
insulin 0.83 IU/kg/day | 588
degludec 50 IU/day | 588
aspart 59 IU/day | 588
oxygen therapy | 588
BiPAP | 588
exercise training | 588
follow-up | 756
HbA1c level 8%–9% | 756
metformin 13.3 mg/kg/day | 756
insulin degludec 76 IU/day | 756
insulin aspart 60 IU/day | 756