79 years old | 0
    male | 0
    lower abdominal pain | 0
    pyrexia | 0
    peri-umbilical pain | -24
    migrated to right lower quadrant pain | 0
    hypertension | 0
    type 2 diabetes mellitus | 0
    hyperlipidaemia | 0
    recent admission for bronchoscopy and biopsy of left bronchial mass | -168
    bronchial carcinoid tumour | -168
    generalized lower abdominal tenderness | 0
    maximal tenderness around periumbilical and right lower quadrant | 0
    abdomen soft | 0
    mild guarding | 0
    active bowel sounds | 0
    no rigidity | 0
    tachycardia (110 beats/min) | 0
    tachypnea (22 times/min) | 0
    mild hypertension (132/78 mmHg) | 0
    pyrexia (38.4 °C) | 0
    normal oxygen saturations (96%) | 0
    no acute confusion | 0
    no neurological deficit | 0
    raised white cell count (16.98 × 103/mm3) | 0
    raised neutrophils | 0
    normal C-reactive protein (0.98 mg/L) | 0
    CT abdomen and pelvis with contrast excluded renal calculi | 0
    dilated tubular structure with mild fat stranding and increased enhancement | 0
    preliminary diagnosis of acute appendicitis | 0
    laparoscopic appendectomy | 24
    intact and mildly erythematous appendix resected | 24
    clear ascitic fluid drained | 24
    acute postoperative deterioration | 24
    increasing oxygen requirements | 24
    consolidation on chest radiograph | 24
    unresolved sepsis concerns | 24
    CT scan review revealed fishbone (1.4 cm) | 24
    microperforation at inferior border of 3rd segment of duodenum | 24
    abscess formation | 24
    fat stranding along right pararenal fascia | 24
    fishbone induced microperforation of duodenum | 24
    retroperitoneal abscess | 24
    exploratory laparotomy | 36
    broad-spectrum intravenous antibiotics (Meropenam) | 36
    laparotomy performed | 36
    retroperitoneal abscess drained | 36
    10 mL pus aspirated | 36
    unable to identify site of perforation and fishbone | 36
    manual pressure applied at presumed site | 36
    area washed out | 36
    retroperitoneal drain inserted | 36
    transferred to intensive care unit | 48
    feeding jejunostomy inserted | 48
    decreasing ventilatory support | 48
    oxygen saturations improved | 48
    chest radiograph resolved | 48
    pain well controlled | 48
    antibiotics converted to oral (levofloxacin) | 48
    retroperitoneal drain removed | 48
    regular oral feeding reintroduced | 48
    discharged after 11 days | 264
    no long-term complications | 264
    jejunostomy tube removed | 264
    pathological examination of appendix showed minimal neutrophils | 48
    excluded acute appendicitis | 48
    abscess cultures isolated intestinal coliforms | 48
    infection from GI source | 48
    initial oxygen desaturation due to pulmonary haemorrhage | 24
    traumatic suctioning during anesthesia | 24
    acute chest radiograph changes | 24
    fishbone attributed to fish soup consumption | -168
    fishbone ingestion not noticed | -168
    <|eot_id|>