56 years old | 0
African American | 0
female | 0
admitted to the Emergency Department | 0
swelling over her left labia | -144
swelling over her left labia developing for six days | -144
swelling opened and begun to drain | -48
temperature was 36.8 ° Celsius | 0
blood pressure was 100/60 mmHg | 0
pulse was 96–100 beats per minute | 0
respiratory rate was 20 breaths per minute | 0
arterial oxygen saturation was 98% | 0
white blood cell count (WBC) was 17.4 × 10^9 per liter | 0
started empirically on vancomycin | 0
started empirically on piperacillin/tazobactam | 0
surgery consult was requested | 0
pelvic CT scan was obtained | 0
cutaneous ulceration over the left labia | 0
air in the subcutaneous fat of the left groin | 0
air in the subcutaneous fat of the left lower abdominal wall | 0
inflammatory fat stranding along the left lateral abdominal wall | 0
LRINEC score was 3 | 0
LRINEC score had the potential to go up to a 7 | 0
decision to perform immediate explorative surgery | 0
explorative surgery of the pelvic and abdominal regions | 2
necrotizing soft tissue infection originating at the left vulva | 2
necrotizing soft tissue infection spreading to the abdominal wall | 2
aggressive debridement | 2
second look exploration surgery | 12
further debridement of the vulvar area | 12
additional pockets of necrosis in the abdominal wall were discovered | 12
additional pockets of necrosis in the abdominal wall were debrided | 12
additional debridement of the genital and abdominal regions | 24
definitive closure of the wound in both areas | 48
stay in the surgical intensive care unit | 0
stay in the surgical intensive care unit was five days long | 120
microbiology samples determined that the offending agents were Clostridium clostridiforme | 24
microbiology samples determined that the offending agents were Bacteroides | 24
Jackson-Pratt drain was placed | 2
Jackson-Pratt drain was removed | 168
patient healed well from the surgery | 168
no complications | 168
proper bowel function | 168
cosmetic outcome was favorable | 168
diagnosis of NF was very challenging | 0
elevated WBC | 0
pelvic CT findings | 0
suspicion of NF | 0
tachycardia | 0
hypotension | 0
despite intravenous fluid resuscitation | 0
despite broad spectrum antibiotic treatment | 0
septic shock | 0
hemodynamic instability | 0
strongest and most valid indicator for emergent surgical exploration | 0
unusual location | 0
lack of associated co-morbidities | 0
lack of risks factors for NF | 0
negative history of initiating trauma | 0
low LRINEC score | 0
cannot be used to eliminate the diagnosis of NF | 0
surgical intervention was performed | 0
prompt surgical debridement | 0
most important and independent prognostic factor | 0
discharged | 168