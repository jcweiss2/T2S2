11 years old | 0  
    girl | 0  
    elective surgery for posterior spinal fusion | -12  
    idiopathic scoliosis | -12  
    anesthesia with propofol | -12  
    estimated blood loss of 1.4 liters | -12  
    received blood products and crystalloid | -12  
    hypotension | -12  
    required packed red blood cells | -12  
    required fresh frozen plasma | -12  
    required cryoprecipitate | -12  
    required platelets | -12  
    vasopressors (phenylephrine and norepinephrine) | -12  
    extubated immediately postoperatively | -12  
    postoperative day 1 | 24  
    disseminated intravascular coagulation | 24  
    liver injury | 24  
    rhabdomyolysis | 24  
    oliguria | 24  
    fluid resuscitation (10 liters) | 24  
    reintubated | 24  
    fluid overload | 24  
    failed response to high-dose diuretics | 24  
    dry weight of 44 kg before surgery | -12  
    weight of 54.6 kg at transfer | 0  
    transferred to tertiary care hospital | 0  
    rhabdomyolysis upon transfer | 0  
    serum creatinine of 4.17 mg/dl | 0  
    creatinine phosphokinase of 17,301 IU/l | 0  
    phosphorus of 9.7 mg/dl | 0  
    uric acid of 10.4 | 0  
    urine myoglobin of 3845 mg/dl | 0  
    acidemic with arterial pH of 7.32 | 0  
    partial pressure of carbon dioxide of 44 mm Hg | 0  
    bicarbonate of 22 mEq/l | 0  
    lactate of 1.7 mmol/l | 0  
    AKI | 0  
    elevated aspartate aminotransferase (3489 IU/l) | 0  
    elevated alanine aminotransferase (2593 IU/l) | 0  
    acute pancreatitis | 0  
    elevated amylase (487 IU/l) | 0  
    elevated lipase (439 IU/l) | 0  
    elevated triglyceride level (135 mg/dl) | 0  
    elevated white blood count | 0  
    DIC | 0  
    elevated protime | 0  
    elevated partial thromboplastin time | 0  
    elevated lactate dehydrogenase (5892 IU/l) | 0  
    elevated d-dimer (>35 mg/dl) | 0  
    low haptoglobin (<10 mg/dl) | 0  
    respiratory failure requiring mechanical ventilation | 0  
    fraction of inspired oxygen of 50% | 0  
    PaO2/fraction of inspired oxygen ratio of 290 | 0  
    not on vasopressors | 0  
    CRRT initiation | 5  
    minimal fluid intake before CRRT | 0  
    fluid overload of 24% at CRRT initiation | 0  
    differential diagnosis of propofol infusion syndrome | 0  
    differential diagnosis of sequelae from intraoperative hypotension | 0  
    met enrollment criteria for SCD trial | 0  
    informed consent provided | 0  
    SCD incorporated into circuit | 7  
    SCD changed every 24 hours | 24  
    stable blood pressure on CRRT and SCD | 24  
    circuit ionized calcium <0.4 mM | 24  
    oxygen requirement stabilized | 24  
    white blood count normalized | 24  
    coagulopathy improved | 24  
    liver injury diminished | 24  
    net fluid volume removal achieved | 24  
    liver enzymes improved | 48  
    pancreatic enzymes improved | 48  
    capillary leak improved | 24  
    net volume removal at 50 ml/h | 48  
    net volume removal at 100 ml/h | 72  
    respiratory function improved | 72  
    extubation | 96  
    temperature spike to 38.4°C | 96  
    elevated white blood count | 120  
    procalcitonin level of 2.64 ng/ml | 120  
    broad spectrum antibiotics started | 120  
    blood cultures negative | 120  
    transition to room air | 168  
    renal function improved | 168  
    completed 7-day SCD treatment | 168  
    no device-related adverse events | 168  
    oliguric at admission | 0  
    nonoliguric with 618 ml/24 h urine output | 240  
    CRRT discontinued | 336  
    transferred to general medical floor | 360  
    discharged home | 480  
    full recovery from liver dysfunction | 480  
    full recovery from lung dysfunction | 480  
    full recovery from kidney dysfunction | 480  
    full recovery from hematologic dysfunction | 480  
    serum creatinine of 0.9 mg/dl at discharge | 480  
    serum creatinine of 0.51 mg/dl at follow-up | 1152  
    