74 years old | 0
male | 0
admitted to the hospital | 0
intermitted fever | -744
progressive back pain | -744
hemoptysis | -744
elevated laboratory values indicating inflammation | -744
ruptured PAU | -744
TEVAR | -744
long-term oral antibiotic therapy | -744
hospitalized | 0
intravenous antibiotic therapy | 0
blood cultures revealed S. aureus | 0
CTA showed gas collections around the aortic stent graft | 0
EI confirmed | 0
infection expanded retrograde right above the celiac trunk | 0
implantation of extra-anatomic ascendobifemoral bypass | 0
counseling with the patient | 0
surgery divided into two stages | 0
minimal sternotomy | 0
AA prepared and clamped tangentially | 0
bypass between AA and left-sided CCA and subclavian artery | 0
aortic arch interrupted distally of the brachiocephalic trunk | 0
ascendobifemoral bypass implanted | 0
proximal end-to-side anastomosis to the AA | 0
anastomosis to both-sided common femoral arteries | 0
left-sided thoracotomy | 0
thoracic abdominal aorta ligated proximal of the celiac trunk | 0
infected stent graft explanted | 0
renal and mesenteric system showed no dysfunctions | 168
inflammation parameters decreased | 168
neurological symptoms did not appear | 168
aspirin and low-molecular-weight heparin therapy established | 168
renal insufficiency with need for dialysis | 720
spondylodiscitis | 720
cholangitis | 720
respiratory insufficiency with prolonged intubation | 720
pneumonia | 720
sepsis | 1440
death | 1440