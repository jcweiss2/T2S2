29 years old | 0
male | 0
admitted to the hospital | 0
biventricular failure | -720
ejection fraction 5-10% | -720
myopericarditis | -720
constrictive physiology | -720
peripherally inserted central catheter (PICC) line placed | -720
discharged on milrinone | -720
fever | -24
chills | -24
septic shock | 0
PICC line removed | 0
IV vancomycin | 0
piperacillin/tazobactam | 0
vasopressor support | 0
Chryseobacterium indologenes grew from PICC line and peripheral blood cultures | 48
antibiotics changed to ciprofloxacin and piperacillin/tazobactam | 48
weaned off vasopressor support | 48
pericardiectomy | 168
completed 14 days of antibiotics | 240
discharged from the hospital | 264
off inotropes | 264
stable vital signs and labs | 264
seen in outpatient cardiology clinic | 744
remains in good health | 744
no evidence of recurrent infection | 744
cardiogenic shock | -720
atrial flutter with rapid ventricular response | -720
radiofrequency ablation | -720
inotrope therapy | -720
home milrinone infusion | -720
follow-up transthoracic echocardiogram | 120
left ventricular EF increased to 50-55% | 120
right ventricular systolic dysfunction improved | 120
furosemide | 0
losartan | 0
metoprolol succinate | 0
milrinone | 0
spironolactone | 0
ciprofloxacin | 48
piperacillin/tazobactam | 0
sacubitril-valsartan | 264
guideline-directed medical therapy for heart failure | 264
no shortness of breath | -24
no chest pain | -24
no redness or drainage around the PICC line | 0
no signs of elevated jugular venous pressure | 0
no lower extremity oedema | 0
bilateral radial and dorsalis pedis pulses were equal and 2+ bilaterally | 0
lungs were clear to auscultation bilaterally | 0
normal work of breathing | 0
fever of 38.7°C | -24
tachycardia with a heart rate in the 110s | -24
blood pressure of 96/57 mmHg | -24
heart was tachycardic, but normal rhythm without any murmurs, rubs, or gallops | -24
Chest X-ray showed no abnormalities | 0
electrocardiogram was significant for sinus tachycardia, normal axis, RSR′ pattern in V1, QRS duration of 90 ms, and non-specific T wave flattening in the inferolateral leads | 0
simultaneous right and left heart catheterization | 120
discordance of the right and left ventricular pressures | 120
diastolic equalization of pressures | 120
supporting the diagnosis of constrictive pericarditis | 120