sixty-nine years old | 0
female | 0
italian | 0
housewife | 0
NLUTD | 0
spondylolisthesis | -1980
surgery for spondylolisthesis | -1980
stress urinary incontinence | -1056
iBC | -1056
recurrent UTIs | -720
problems during monthly iBC change | -720
abdominal cross-sectional imaging | 0
ultrasound | 0
computed tomography | 0
bladder stone | 0
videourodynamic study | 0
defunctionalized bladder | 0
uterus-sparing simple cystectomy | 0
uretero-ileal-cutaneous diversion | 0
antibiotic prophylaxis | 0
Cefazolin | 0
operative time | 0
septic | 72
severe lumbar pain | 72
abdominal fluid cultures | 72
Escherichia coli | 72
Pseudomonas aeruginosa | 72
Candida glabrata | 72
pancreatic oedema | 72
conservative approach | 72
septic shock | 432
Enterococcus faecium | 432
Acinetobacter spp | 432
urgent exploratory laparotomy | 432
acute necrotizing hemorrhagic pancreatitis | 432
medical therapy | 432
abdominopelvic washing | 432
septic episodes | 432
discharged | 141*24
well-functioning urinary diversion | 141*24+2*365*24
no significant conditions in urinary tract | 141*24+2*365*24