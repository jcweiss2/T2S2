62 years old | 0
male | 0
admitted to the hospital | 0
progressive debilitating fatigue | -72
diffuse skin lesions | -72
generalized lymphadenopathy | -72
anemic | -72
blasts in peripheral blood | -72
extensive axillary lymphadenopathy | -72
mediastinal lymphadenopathy | -72
inguinal lymphadenopathy | -72
splenomegaly | -72
monocytic precursors expressing CD56 and CD123 | -72
bone marrow biopsy | -72
bone marrow aspiration | -72
blasts in bone marrow | -72
CD7 positive | -72
CD33 positive | -72
CD38 positive | -72
CD56 positive | -72
CD71 positive | -72
CD117 positive | -72
CD123 positive | -72
HLA-DR positive | -72
CD3 negative | -72
CD4 negative | -72
CD10 negative | -72
CD19 negative | -72
CD34 negative | -72
MPO negative | -72
TdT negative | -72
skin biopsy | -72
fine needle aspiration of inguinal nodes | -72
tagraxofusp treatment | 0
recurrent scalp lesion | 144
biopsy of recurrent scalp lesion | 144
Hyper-CVAD treatment | 168
neutropenic fever | 192
progressive hypoxia | 192
hospitalized | 192
intensive care unit (ICU) level of care | 192
broad spectrum antibiotics | 192
steroid course | 192
drug-induced pneumonitis | 192
cyclophosphamide | 192
cerebrospinal fluid (CSF) analysis | 192
blasts in CSF | 192
intrathecal (IT) methotrexate therapy | 192
CD34+ allogenic stem cell transplant | 240
fludarabine | 240
melphalan | 240
engraftment syndrome | 264
Staphylococcal epidermidis bacteremia | 264
Clostridium difficile infection | 264
angioedema | 264
generalized exanthematous pustulosis | 264
ICU level of care | 264
bone marrow repeated | 288
recurrent BPDCN | 288
47.5% blasts in bone marrow | 288
CSF positive for disease | 288
vyxeos treatment | 312
IT methotrexate continued | 312
bone marrow aspirate | 336
complete response to vyxeos | 336
no evidence of BPDCN | 336
neutropenic fever | 360
pseudomonas infection | 360
sepsis | 360
overwhelming infection | 360
death | 360