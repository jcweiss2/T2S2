54 years old | 0
male | 0
decompensated nonalcoholic steatohepatitis cirrhosis | -672
OLT | -672
side-to-side cavoplasty | -672
duct-to-duct biliary anastomosis | -672
end-to-end portal vein anastomosis | -672
end-to-end common HA anastomosis | -672
discharged home | -504
physical therapy | -504
syncope | -24
fall | -24
trimalleolar left ankle fracture | -24
ibuprofen | -168
arthralgias | -168
dark stools | 0
vomiting fresh blood with clots | 0
5 g drop in hemoglobin | 0
intubated | 0
urgent upper endoscopy | 0
hemorrhagic shock | 0
gastrointestinal hemorrhage | 0
resuscitated with blood products | 0
cratered 2–3 cm ulcer in the proximal duodenum | 0
large vessel visible | 0
endoscopic therapy with 1.2 mL of epinephrine injection | 0
endoscopic therapy with 2 endoclips | 0
endoscopic therapy with 1 minute of bipolar electrocautery | 0
antral biopsies not obtained | 0
Stool Helicobacter pylori testing recommended | 0
mesenteric angiogram | 12
possible embolization | 12
luminal narrowing and irregularity of the proper HA | 12
nonfilling of the GDA | 12
aspartate aminotransferase of 2,686 U/L | 12
alanine aminotransferase of 3,406 U/L | 12
ischemic hepatitis | 12
computed tomography angiogram | 24
severe proper HA stenosis | 24
moderate common HA stenosis | 24
GDA occlusion | 24
multifocal hepatic infarcts | 24
thickening in the first part of the duodenum | 24
surgical intervention | 24
exploratory laparotomy | 48
duodenum adherent to the donor HA | 48
full-thickness ulceration of the superior aspect of the duodenum | 48
HA pseudoaneurysm | 48
proximal and distal control gained | 48
aneurysmal segment resected | 48
new end-to-end anastomosis created | 48
ultrasound demonstrated excellent flow | 48
Graham patch sutured onto the duodenum | 48
right upper quadrant drain placed | 48
abdomen closed | 48
transferred to the intensive care unit | 48
intubated | 48
stable condition | 48
perioperative antibiotics | 48
abdominal fluid cultures positive for Streptococcus mitis group | 48
abdominal fluid cultures positive for Haemophilus influenzae | 48
extubated | 72
open reduction and internal fixation of the left trimalleolar ankle fracture | 96
liver functions normalized | 96
repeat liver ultrasound demonstrated normal flow through the transplant HA | 96
discharged to a subacute rehab facility | 312
medically stable | 312