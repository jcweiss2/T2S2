nursing student reported | 0
outpatient department | 0
fever | -48
vesicular lesions | -48
face | -48
chest | -48
back | -48
whole body | -48
varicella infection | 0
denied being in contact with a chicken pox infected case | 0
attending a patient with HZ infection | -336
not immune to varicella infection | 0
neither vaccinated nor had been infected with varicella virus previously | 0
fluid from the blisters | 0
sent for serological examination | 0
confirmed the diagnosis of VZV infection | 48
two staff nurses | 48
medicine resident doctor | 48
similar history | 48
clinical manifestations | 48
four more health care workers | 120
fever | 120
vesicular lesions | 120
started on treatment | 120
granted leave from duty | 120
reported to infection control committee | 120
reported to administration | 120
investigation of the outbreak | 120
probable index case | -672
60-year-old male | -672
admitted | -672
road side accident | -672
blunt trauma chest | -672
rib fractures | -672
right intercostal drain | -672
right lower zone pneumonia | -672
renal failure | -672
left ventricular dysfunction | -672
septic shock | -576
despite antibiotic cover | -576
resuscitative measures | -576
skin lesions | -336
right L2, 3, 4 dermatome | -336
skin consultation | -336
lesions identified as localized HZ | -336
started on tab acyclovir | -336
T-bact ointment dressings | -336
succumbed to septic shock | -240
multiorgan failure | -240
expired | -240
eight HCWs infected | 336
directly or indirectly involved in care of the index case | 336
rest of the susceptible staff | 336
vaccinated with chickenpox vaccine | 336
old and new patients | 336
screened and tracked | 336
did not develop any such lesions | 720
no new VZV infection | 720
among HCWs | 720
among patients | 720
varicella is highly contagious | 0
average incubation period | 0
 Persons with varicella are considered infectious | 0
from 1 to 2 days before the rash appears | 0
until all lesions are crusted over | 0
outbreak of varicella | 0
five or more cases | 0
specific setting | 0
epidemiologically linked | 0
surveillance | 0
through two full incubation periods | 0
after the rash onset | 0
last identified case-patient | 0
reactivation of latent VZV | 0
results in HZ infection | 0
shingles | 0
patients with zoster | 0
contagious to those who have no immunity to VZV | 0
route of transmission | 0
via direct contact | 0
exposure to dressings | 0
clothing soiled with blister fluid | 0
current guidelines | 0
prevention of varicella spread | 0
from a HZ patient | 0
standard infection-control precautions | 0
covering of HZ lesions | 0
means of preventing nosocomial spread | 0
do not recommend the isolation | 0
all affected patients | 0
airborne transmission | 0
may occur | 0
varicella | 0
zoster | 0
strategies for managing zoster patients | 0
same precautions | 0
airborne transmission | 0
varicella patients | 0
reduce the risk for transmission | 0
vaccination for chickenpox | 0
not included in National Immunization schedule | 0
recommended by Indian Academy of Pediatrics | 0
chickenpox in adults | 0
more severe than in children | 0
better to get the children vaccinated | 0
unvaccinated VZV exposed healthcare personnel | 0
without evidence of VZV immunity | 0
receive postexposure vaccination | 0
as soon as possible | 0
vaccination within 3–5 days | 0
of exposure to rash | 0
modify the disease | 0
if infection occurred | 0
vaccination 6 or more days | 0
after exposure | 0
still indicated | 0
induces protection | 0
against subsequent exposures | 0
second dose | 0
given 4–6 weeks | 0
after the first dose | 0
unvaccinated VZV-susceptible healthcare personnel | 0
at risk for severe disease | 0
varicella vaccination | 0
contraindicated | 0
e.g. pregnant healthcare personnel | 0
varicella-zoster immune globulin | 0
after exposure | 0
breach in infection control precautions | 0
caused varicella outbreak | 0
in our ICU | 0
made certain changes | 0
in our hospital policy | 0
prevent a future outbreak | 0
healthcare personnel | 0
alerted to the risks | 0
possible infection | 0
offered 2 doses | 0
of varicella vaccine | 0
when they begin employment | 0
stringent airborne | 0
contact precautions | 0
ensured | 0
not only in patients | 0
suffering from varicella | 0
but also in patients | 0
with HZ infection | 0
in future | 0