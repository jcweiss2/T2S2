76 years old | 0
renal transplant woman | 0
admitted to the Intensive Care Unit (ICU) | 0
coma | 0
respiratory distress | 0
methylprednisolone | 0
tacrolimus | 0
mycophenolate mofetil | 0
candesartan | 0
arterial hypertension | 0
serum creatinine concentration 1.70 mg/dl | -432
estimated glomerular filtration rate (GFR) 28 ml/min/1.73 m2 | -432
Hepatitis B virus (HBV) reactivation | -12960
109 DNA copies/ml | -12960
no specific treatment | -12960
liver tests within normal range | -12960
progressive dyspnea | -288
chest X-ray | -288
lung computed tomography (CT) | -288
bilateral lung infiltrates | -288
cytomegalovirus (CMV) polymerase chain reaction (PCR) in plasma 3130 copies/ml | -288
culture of the bronchoalveolar lavage | -288
diagnosis of CMV pneumonia | -288
intravenous sodium ganciclovir | -288
initial daily dose of 200 mg | -288
increased to 400 mg (4.2 mg/kg) | -264
CMV PCR became rapidly negative | -264
white blood cell count 5080/mm3 | -288
nadir at 3430/mm3 | -264
renal function deteriorated | 0
creatinine 2.67 mg/dl | 0
estimated GFR declining from 26 to 17 ml/min/1.73 m2 | 0
hip fracture | 288
orthopedic surgery | 288
epidural anesthesia | 288
altered consciousness | 288
respiratory distress | 288
arterial blood gas analysis | 288
pH 6.79 | 288
pCO2 54 mm Hg | 288
bicarbonate 8 mmol/l | 288
lactate 20 mmol/l | 288
intubated for mechanical ventilation | 288
intravenous 8.4% sodium bicarbonate | 288
thiamine supplementation | 288
continuous venovenous hemofiltration | 288
arterial pH rose progressively up to 7.31 | 294
central venous oxygen saturation (ScvO2) 61.5% | 294
echocardiography showed well preserved left ventricular function | 294
no evidence for septic shock | 294
no evidence for hemorrhagic shock | 294
arterial lactate (L) 27 mmol/l | 294
pyruvate (P) 0.6 mmol/l | 294
L/P molar ratio 45 | 294
hypoglycemia | 294
administration of dextrose 30% | 294
impaired glucose utilization | 294
biological signs of ketogenesis | 294
high urinary excretion of 3-hydroxybutyrate 256.2 mmol/mol creatinine | 294
high urinary excretion of dicarboxylic acids | 294
ganciclovir therapy discontinued | 288
11-day course | -288
rhabdomyolysis | 288
vasoplegia | 288
blood cultures sterile | 288
abdominal CT showed no sign of bowel ischemia | 288
hyperlactatemia | 288
liver tests moderately disturbed | 288
ammonia level 109 μg/dl | 288
severely encephalopathic | 288
normal brain CT | 288
fatality | 336
persisting hyperlactatemia (>25 mmol/l) | 336
circulatory failure | 336
progressive increase of vasopressors | 336
autopsy not accepted | 336
