57 years old | 0
male | 0
lepromatous leprosy | -60
skin biopsy | -60
treatment with rifampicin/clofazimine/dapsone | -60
admitted to the hospital | 0
abdominal distension | 0
constipation | 0
vomiting | 0
10-kg weight loss | 0
peripheral lymphadenopathy | 0
distended abdomen | 0
positive shifting dullness | 0
computed tomography scan of abdomen | 0
mural thickening of terminal ileum | 0
enlarged mesenteric lymph nodes | 0
mesenteric fat stranding | 0
intra-abdominal free fluid | 0
abdominal paracentesis | 0
atypically large lymphocytes | 0
flow cytometry | 0
abnormal CD4/CD8 double-negative T-cell population | 0
cervical lymph node biopsy | 0
high-grade peripheral T-cell lymphoma | 0
bone marrow examination | 0
no involvement of T-cell NHL | 0
stage IV lymphoma | 0
dexamethasone | 0
tumor-lysis syndrome precautions | 0
deteriorated clinically | 24
transferred to medical ICU | 24
severe sepsis | 24
antibiotics | 24
antifungals | 24
ICU care | 24-168
recovered | 168
transferred to national cancer center | 168
EPOCH chemotherapy protocol | 168
CNS prophylaxis | 168
intrathecal methotrexate | 168
febrile neutropenia episodes | 336
recurrent bacteremia | 336
generalized weakness | 336
no sensory changes | 336
no clear fatigability | 336
decreased power in proximal and distal muscles | 336
normal distal latencies | 336
normal compound muscle action potential | 336
normal conduction velocities | 336
normal F waves | 336
normal sensory nerve studies | 336
needle electromyogram | 336
poor recruitment effects | 336
repetitive nerve stimulation | 336
significant incremental response | 336
presynaptic neuromuscular junction disorder | 336
LEMS | 336
intravenous immunoglobulins | 336
significant improvement of motor function | 360
ambulate | 360
planned for consolidation by autologous bone marrow transplant | 360
recurrent bacteremia and sepsis | 720
re-admitted to medical ICU | 720
severe sepsis and multiorgan failure | 720
passed away | 1440