20 years old | 0
    male | 0
    diagnosed with schizophrenia | 0
    diagnosed with cannabis use disorder | 0
    diagnosed with social anxiety disorder | 0
    delusional belief | 0
    fecal odour | 0
    risperidone | -17520
    paliperidone palmitate | -17520
    quetiapine | -17520
    CGI-S score 5 | -17520
    weight gain 35 kg | -17520
    clozapine initiation | -4320
    CGI-S score 3 | -4320
    cannabis use disorder remission | -4320
    weight gain 10 kg | -4320
    sertraline initiation | -4320
    clozapine dose increase | -240
    muscular pain | -240
    CK level 7,499 U/L | -240
    weight training | -240
    transferred to medical facility | 0
    clozapine stopped | 0
    benztropine introduction | 0
    aggressive fluid therapy | 0
    clozapine levels normal | 0
    recreational drug negative | 0
    myocarditis ruled out | 0
    NMS ruled out | 0
    denies performance enhancement drugs | 0
    overweight | 0
    CK peak 45,564 U/L | 72
    CK normalized | 336
    discharged | 336
    sertraline discontinued | 336
    aripiprazole | 336
    lorazepam | 336
    CGI-S score 6 | 336
    visual hallucinations | 336
    auditory hallucinations | 336
    clozapine rechallenge | 2976
    CK monitoring | 2976
    clozapine reinitiation | 2976
    CK level 2,218 U/L | 2976
    weight training | 2976
    clozapine continued | 2976
    CK normalized | 2976
    weight training | 2976
    CK level 4,734 U/L | 2976
    CK normalized | 2976
    CGI-S score 3 | 2976
    