66 years old | 0
male | 0
diabetes mellitus type 2 | 0
hypertension | 0
dyslipidemia | 0
admitted to the hospital | 0
dry cough | -168
mild shortness of breath | -168
fever | -168
discharged home | -168
reverse transcription–polymerase chain reaction (RT-PCR) test | -168
SARS-CoV-2 positive | -168
returned to the hospital | -168
worsening shortness of breath | -168
transferred to the institution | -168
admitted to the intensive care unit | 0
hydroxychloroquine treatment | 0
azithromycin treatment | 0
intravenous (IV) ceftriaxone treatment | 0
respiratory distress | 96
severe hypoxia | 96
oxygen saturation 40% | 96
hemodynamically unstable | 96
blood pressure 50/31 mm Hg | 96
intubated | 96
resuscitated with 2 liters of IV fluid boluses | 96
norepinephrine infusion | 96
vasopressin infusion | 96
epinephrine infusion | 96
point-of-care cardiac ultrasonography | 96
severely reduced LVEF | 96
dobutamine treatment | 96
arterial blood gas | 96
pH 7.17 | 96
PaCO2 48 | 96
PaO2 69 | 96
bicarbonate 19 mmol/L | 96
FiO2 100% | 96
PaO2/FiO2 ratio 69 | 96
chest X-ray | 96
interval worsening of patchy and confluent opacities | 96
electrocardiogram (ECG) | 96
sinus tachycardia | 96
low voltage complexes | 96
nonspecific T-wave abnormalities | 96
troponin T 0.39 ng/mL | 96
NT-proBNP 798 pg/mL | 96
transthoracic echocardiography | 120
normal LV size | 120
severe LV dysfunction | 120
estimated LVEF 32% | 120
global LV hypokinesia | 120
ferritin 100586 ng/mL | 120
lactate dehydrogenase (LD) >25000 U/L | 120
D-dimer 6.99 µg/mL | 120
C-reactive protein (CRP) 278.4 mg/L | 120
convalescent plasma administration | 120
convalescent plasma administration | 144
norepinephrine infusion discontinued | 120
vasopressin infusion discontinued | 120
epinephrine infusion discontinued | 120
dobutamine infusion deescalated | 120
mechanical ventilation | 120
antibiotics (IV vancomycin and cefepime) | 120
IV diuretics | 120
cardiogenic shock improved | 192
dobutamine infusion discontinued | 192
troponin T 0.05 ng/mL | 192
NT-proBNP 26 pg/mL | 192
ferritin 4320 ng/mL | 192
CRP 69.7 mg/L | 192
D-dimer 2.38 µg/mL | 192
LD 427 U/L | 192
transthoracic echocardiography | 240
improved LVEF (60% to 65%) | 240
normal LV systolic function | 240
no wall motion abnormalities | 240
extubated | 360
COVID-19 RT-PCR test negative | 456
discharged home | 504