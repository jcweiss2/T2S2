83 years old | 0
    woman | 0
    insulin-dependent diabetes mellitus | -3
    hypertension | -3
    hyperlipidemia | -3
    diastolic heart failure | -3
    diabetic gastroparesis | -3
    chronic kidney disease | -3
    nausea | -72
    substernal epigastric abdominal discomfort | -72
    belching | -72
    poor oral intake | -72
    mild right upper quadrant tenderness | 0
    aperistalsis of the esophageal body | 0
    elevated LES pressure | 0
    type I achalasia | 0
    decreased motility of the esophagus | 0
    underwent esophagogastroduodenoscopy | 0
    botulinum toxin injections targeting LES | 0
    discharged | 0
    right shoulder pain | 504
    given NSAIDS | 504
    symptoms persisted | 504
    referred to pain specialist | 504
    right shoulder intra2-articular steroid injections | 504
    prescribed NSAIDS | 504
    symptoms continued | 504
    presented to emergency department | 528
    white blood cell count 30.7 K/μL | 528
    computed tomography scan of abdomen | 528
    5.8 cm x 6.9 cm x 2.3 cm fluid collection | 528
    abscess near diaphragm | 528
    started on vancomycin | 528
    started on piperacillin/tazobactam | 528
    abscess drained | 528
    fluid cultures grew Streptococcus intermedius | 528
    vancomycin trough after third dose 32 μg/ml | 528
    vancomycin discontinued | 528
    piperacillin/tazobactam discontinued | 528
    started on ampicillin/sulbactam | 528
    leukocytosis improved | 528
    repeat abdominal CT | 528
    interval decrease in abscess size | 528
    generalized edema | 528
    acute kidney injury | 528
    hemodialysis initiated | 528
    unresponsive during hemodialysis | 528
    endotracheal intubation | 528
    admitted to medical intensive care unit | 528
    septic shock | 528
    vasopressor support | 528
    antibiotics escalated to meropenem | 528
    antibiotics escalated to vancomycin | 528
    ischemic hepatopathy | 528
    large left pleural effusion | 528
    chest tube placement | 528
    atrial fibrillation with rapid ventricular response | 528
    placed on comfort care measures | 840
    died | 840
