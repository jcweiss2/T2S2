23 years old | 0
female | 0
sore throat | -72
nausea | -72
subjective fever | -72
chills | -72
given oral antibiotics | -24
febrile | 0
tachycardic | 0
hypotensive | 0
leukocyte count of 17.87 k/ul | 0
neutrophil count of 86.8% | 0
elevated creatinine of 3.6 mg/dL | 0
sepsis | 0
acute kidney injury | 0
empiric antibiotics | 0
rapid crystalloid infusion | 0
hypotensive | 0
admitted to the intensive care unit | 0
fulminant septic shock | 0
Streptococcus anginosus isolated from blood cultures | 0
F. necrophorum isolated from blood cultures | 0
scattered bilateral nodular opacities throughout the lung | 0
septic emboli | 0
small bilateral pleural effusions | 0
adjacent consolidations | 0
piperacillin/tazobactam | 0
metronidazole | 0
Lemierre's syndrome suspected | 0
internal jugular vein thrombosis ruled out | 0
decrease in the size of the bilateral nodular opacities | 240
new areas of cavitation | 240
increased moderate left pleural effusion | 240
near complete atelectasis of the left lower lobe | 240
Left sided chest tube placed | 240
parapneumonic effusion | 240
F. necrophorum sensitive to augmentin | 240
F. necrophorum sensitive to clindamycin | 240
F. necrophorum sensitive to imipenem | 240
F. necrophorum resistant to metronidazole | 240
Streptococcus anginosus pansensitive to penicillin | 240
Streptococcus anginosus pansensitive to ceftriaxone | 240
Streptococcus anginosus pansensitive to clindamycin | 240
Streptococcus anginosus pansensitive to vancomycin | 240
Streptococcus anginosus pansensitive to levofloxacin | 240
Streptococcus anginosus pansensitive to erythromycin | 240
antibiotics switched to piperacillin/tazobactam and clindamycin | 240
diagnosed with Lemierre's syndrome | 240
pulmonary septic emboli | 240
discharged home | 432
ceftriaxone | 432
clindamycin | 432
good recovery | 432