79 years old | 0
female | 0
admitted to the hospital | 0
fever | -120
malaise | -120
anorexia | -120
confusion | -72
unconsciousness | -72
diabetes | -16560
hypertension | -16560
atrial fibrillation | -16560
cholecystectomy | -16560
appendectomy | -16560
pyrexia | 0
noninvasive mechanical ventilation | 0
tachycardia | 0
decreased breath sounds | 0
soft abdomen | 0
no peripheral edema | 0
increased procalcitonin level | 0
high white blood cell count | 0
anemia | 0
low platelet cell count | 0
elevated N-terminal pro-B-type natriuretic peptide levels | 0
liver abscess | -120
hepatic venous gas | 0
gas bubbles in the hepatic vein | 0
gas bubbles in the inferior vena cava | 0
gas bubbles in the right atrium | 0
ruptured liver abscess | 0
Klebsiella pneumoniae infection | 0
imipenem and cilastatin treatment | 0
cefoperazone sulbactam treatment | 120
improvement of infection index | 168
no further gas in the hepatic vein | 48
small liquefaction zone in the abscess area | 48
abscess shrinkage | 168
abscess disappearance | 984
discharged from the hospital | 984