71 years old | 0
female | 0
metastatic renal cell carcinoma (mixed papillary and clear cell type) | 0
retroperitoneal lymph node metastasis | 0
right ovarian metastasis | 0
liver metastasis | 0
first-line doublet immunotherapy with ipilimumab and nivolumab | 0
maintenance single-agent nivolumab | 0
immune-related primary hypoadrenalism | 0
immune-related hypopituitarism | 0
secondary hypoadrenalism | 0
hypothyroidism | 0
exogenous hydrocortisone | 0
fludrocortisone | 0
thyroxine replacement | 0
short synacthen test | 0
MRI pituitary | 0
disease progression | 0
second-line sunitinib | 0
admitted to the hospital with presumed sepsis | 336
fever | 336
hypotension | 336
tachycardia | 336
broad-spectrum antibiotics | 336
intravenous stress dose steroids | 336
inotropes in the intensive care unit | 336
septic screen | 336
recovered fully | 336
discharged from the hospital | 336
steroid replacement adjusted | 336
sunitinib restarted | 336
re-presented with same symptoms | 432
managed for sepsis | 432
intravenous stress dose steroids | 432
inotropes in ICU | 432
transthoracic echocardiogram | 432
baseline steroid dose reviewed | 432
recommenced on reduced dose of sunitinib | 432
re-presented with same symptoms | 480
ICU admission | 480
stress dose steroids | 480
inotropes | 480
broad-spectrum antibiotics | 480
septic screen negative | 480
tunnelled venous access catheter removed | 480
baseline steroid dose revised | 480
elective admission for trial of sunitinib | 576
sunitinib administration | 576
profoundly hypotensive | 576
tachycardic | 576
intravenous fluid replacement | 576
intravenous steroids | 576
inotropes | 576
haemodynamic parameters normalized | 600
transitioned back to oral steroids | 600
sunitinib therapy permanently discontinued | 600
no fevers recorded | 0
subjective chills | 0
greater than 1° temperature rise | 576
adrenal crisis | 576
adrenal crisis with each rechallenge of sunitinib | 432 | 480 | 576
residual adrenal function insufficient | 0
negative adrenal tissue antibody | 0
negative septic screens | 336 | 432 | 480 | 576
sunitinib-induced adrenal crisis | 336 | 432 | 480 | 576
hypoadrenalism | 0
no conflicts of interest | 0
no funding received | 0
