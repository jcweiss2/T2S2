19 years old | 0
male | 0
admitted to the hospital | 0
paraquat ingestion | -2
nausea | -2
vomiting | -2
Glasgow Coma scale normal | 0
vital signs normal | 0
blood pressure 120/80 mmHg | 0
pulse rate 90/min | 0
respiratory rate 18/min | 0
temperature 37°C | 0
O2 saturation 95% | 0
hypothyroidism | -672
levothyroxine tablets | -672
nasogastric tube | 0
gastrointestinal washing | 0
activated charcoal | 0
dithionite test positive | 0
hemodialysis | 0
N-acetylcysteine administration | 0
Vitamin C infusion | 0
Vitamin E injection | 0
methylprednisolone IV | 0
pantoprazole ampule | 0
silymarin | 0
cervical pain | 504
breathing difficulty | 504
cervical emphysema | 504
chest X-ray | 504
lateral neck graphy | 504
bilateral pneumothorax | 504
pneumomediastinum | 504
bilateral chest tube | 504
fever | 504
pulmonary infection | 504
sepsis | 504
broad-spectrum antibiotic | 504
ALT abnormal | 288
ALT normal | 552
AST normal | 0
AST abnormal | 648
BUN abnormal | 96
BUN fluctuation | 504
creatinine abnormal | 72
creatinine increased | 264
Hb less than normal | 0
anemia | 0
platelet level abnormal | 504
INR abnormal | 648
death | 648
subcutaneous emphysema | 504
pneumothorax | 504
pneumomediastinum severe | 648