18 years old | 0
male | 0
history of intravenous drug use | -168
history of attention deficit/hyperactivity disorder | -168
fever | -168
chills | -168
shortness of breath | -168
non-smoker | -168
no alcohol consumption | -168
fentanyl abuse | -168
dextroamphetamine/amphetamine | -168
admitted to the hospital | 0
fever | -72
chills | -72
shortness of breath | -72
temperature 102.7°F | 0
blood pressure 102/56 mmHg | 0
pulse 136 beats per minute | 0
respiratory rate 38 breaths per minute | 0
oxygen saturation 94% | 0
bilateral rhonchi | 0
tachycardia | 0
no murmur, rub or gallop | 0
white blood cell count 12,200/mm3 | 0
hemoglobin 10.9 g/dL | 0
platelet count 85,000/mm3 | 0
ESR 60 mm/hr | 0
hyponatremia | 0
sodium 124 mmol/L | 0
creatinine level 2.8 mg/dL | 0
BUN 98 mg/dL | 0
NT-proBNP 1028 pg/mL | 0
ECG sinus tachycardia | 0
chest radiograph bilateral lower lobe infiltrates | 0
small pleural effusions | 0
IV fluids | 0
levofloxacin | 0
community acquired pneumonia | 0
septic shock | 0
acute respiratory failure | 0
pressor support | 0
mechanical ventilation | 0
blood cultures gram-positive cocci | 0
vancomycin | 0
tricuspid valve vegetation | 0
tricuspid regurgitation | 0
cardiothoracic surgery | 0
transesophageal echocardiogram | 0
patent foramen ovale | 0
shunt | 0
CT chest multiple cavitary peripheral lung nodules | 0
septic emboli | 0
non-oliguric AKI | 0
renal replacement therapy | 0
acute tubular necrosis | 0
methicillin sensitive Staphylococcus aureus | 0
oxacillin | 0
improved on supportive and antimicrobial therapy | 0
weaned off pressors | 0
successfully extubated | 0
renal function recovered | 0
bilateral nontender purpuric papules | 12
bullous lesions | 12
HIV antibody negative | 12
hepatitis B serology negative | 12
p-ANCA negative | 12
c-ANCA negative | 12
cryoglobulin negative | 12
rheumatoid factor negative | 12
ANA weakly positive | 12
anti-ds DNA antibody negative | 12
Complement C3 low | 12
Complement C4 low | 12
anti-HCV antibody positive | 12
HCV viral load 4.16 × 10^5 IU/mL | 12
aspirated fluid from bullous lesions | 12
no bacteria | 12
no organisms seen on gram staining | 12
punch biopsies from bullous skin lesions | 12
perivascular neutrophil infiltration | 12
fibrinoid necrosis of small vessels | 12
leukocytoclastic vasculitis | 12
vancomycin | 12
resolution of skin lesions | 12
tricuspid valve replacement surgery | 24
no perioperative complications | 24
no recurrence of skin lesions | 30