22 years old | 0
male | 0
admitted to the hospital | 0
pain in the left upper abdomen | -48
shortness of breath | -48
past history of repeated episodes of mild to moderate breathlessness | -672
symptomatic treatment | -672
chest radiograph | -48
air fluid level in the left hemithorax | -48
hydropneumothorax | -48
left-sided intercostal drain (ICD) inserted | -48
serosanguinous fluid drained | -48
second ICD inserted | -24
fluid stained with blood drained | -24
temporary relief of respiratory symptoms | -24
low-grade fever | -24
pleuritic chest pain | -24
referred to hospital | -24
unable to pass stool or flatus | -48
non-bilious vomiting | -48
febrile | 0
hemodynamically stable | 0
two left ICDs in the left hemithorax | 0
turbid, foul-smelling contents drained | 0
decreased air entry on the left side of the lung | 0
abdominal viscera and fluid in the left hemithorax | 0
abdominal tenderness | 0
guarding and rigidity | 0
respiratory embarrassment | 0
absent bowel sounds | 0
pulse rate 122 per min | 0
blood pressure 90 mm Hg systolic | 0
respiratory rate 34–36 per min | 0
pulse oximetry saturation 92–94% | 0
blood investigations unremarkable | 0
mild hypoxemia | 0
mild metabolic acidosis | 0
chest radiograph with air-fluid level | 0
emergency exploratory laparotomy | 0
general anesthesia induced | 0
crash induction performed | 0
intubated with cuffed oral endotracheal tube | 0
maintained on oxygen, nitrous oxide and isoflurane | 0
intravenous fluids infused | 0
20×10 sq cm defect in the posterolateral part of the left dome of the diaphragm | 0
stomach, splenic flexure of the colon and spleen herniated into the left side of the chest | 0
no peritoneal sac over the stomach | 0
ICDs traumatized the spleen and stomach | 0
ICDs removed | 0
splenectomy done | 0
hernial contents reduced | 0
perforation in the stomach closed | 0
ICD placed in the pleural cavity | 0
diaphragmatic defect repaired | 0
transfusion of two units of packed red blood cells | 0
shifted to intensive care unit | 0
respiratory and hemodynamic support | 0
reversal of neuromuscular blockade not done | 0
mild pleural effusion in the left hemithorax | 24
lung re-expanded on serial chest radiographs | 72
extubated on the fifth postoperative day | 120
hemodynamically stable | 120
chest expansion techniques and physiotherapy | 120
transferred to general ward on the seventh postoperative day | 168
recovered without further complications | 168