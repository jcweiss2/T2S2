63 years old | 0  
    woman | 0  
    transient ischemic attack | -6720  
    reflux | -6720  
    hypertension | -6720  
    hyperlipidemia | -6720  
    laparoscopic sleeve gastrectomy | -6720  
    vitamin supplements | -6720  
    weight loss | -6720  
    weight gain | -6720  
    GERD symptoms | -72  
    large hiatal hernia | -72  
    laparoscopic hand-assisted hiatal hernia repair | -72  
    conversion of sleeve gastrectomy to Roux-en-Y gastric bypass | -72  
    adhesive disease | -72  
    uncomplicated procedure | -72  
    inpatient postoperative course | -72  
    discharged home | -72  
    POD 4 | -72  
    outpatient bariatric institute follow-up | -72  
    POD 8 | -72  
    shortness of breath | 432  
    left lower leg pain | 432  
    swelling | 432  
    hypotensive | 432  
    unresponsive | 432  
    cardiopulmonary arrest | 432  
    cardiopulmonary resuscitation | 432  
    return of spontaneous circulation | 432  
    intubated | 432  
    rapid sequence intubation | 432  
    admitted to ICU | 432  
    acidotic | 432  
    pH 7.19 | 432  
    bicarbonate 10 | 432  
    lactic acid 17 | 432  
    base excess −16.4 | 432  
    acute hypoxic respiratory failure | 432  
    renal failure | 432  
    CT imaging | 432  
    pulmonary embolism protocol | 432  
    enlarged left common iliac veins | 432  
    enlarged external iliac veins | 432  
    enlarged common femoral veins | 432  
    edema of left thigh | 432  
    ICU transfer | 432  
    general surgery consultation | 432  
    left leg swelling | 432  
    purple discoloration | 432  
    cold to touch | 432  
    therapeutic anticoagulation | 432  
    vascular surgery consultation | 432  
    PCD concern | 432  
    clinical status not improving | 432  
    diagnostic laparoscopy | 432  
    lower-extremity venogram | 432  
    OR on anticoagulation | 432  
    pink viable bowel | 432  
    no abnormalities | 432  
    venogram via left popliteal vein | 432  
    8-French catheter | 432  
    extensive acute left iliac venous thrombosis | 432  
    femoral venous thrombosis | 432  
    iliac confluence to distal femoral vein | 432  
    thrombectomy | 432  
    clot retrieval system | 432  
    thrombus removal | 432  
    completion venogram | 432  
    clinical status deterioration | 432  
    multisystem organ failure | 432  
    shock liver | 432  
    respiratory failure | 432  
    disseminated intravascular coagulation | 432  
    increasing vasopressor support | 432  
    significant acidosis | 432  
    continuous renal replacement therapy | 432  
    worsening renal failure | 432  
    POD 1 | 504  
    tense left lower extremity | 504  
    bullous formation | 504  
    mottled digits | 504  
    no pulses | 504  
    no Doppler signals | 504  
    compartment syndrome suspicion | 504  
    calf fasciotomy | 504  
    viable muscle | 504  
    thigh fasciotomy | 504  
    copious brown fluid | 504  
    pale muscle | 504  
    tissue death | 504  
    transferred back to ICU | 504  
    cardiopulmonary arrest recurrence | 504  
    resuscitation attempt | 504  
    death | 504  
    multisystem organ failure | 504  
    reperfusion injury | 504  
    VTE complication | 504  
    phlegmasia cerulea dolens | 504  
    postoperative complications | 504  
    reoperation | 504  
    ICU admission | 504  
    readmission | 504  
    end-organ dysfunction | 504  
    mortality | 504  
    therapeutic anticoagulation | 504  
    mechanical thrombectomy | 504  
    amputation | 504  
    fatal reperfusion injury | 504  
    underdiagnosed VTE | 504  
    increased VTE risk | 504  
    early recognition | 504  
    intervention | 504  
    limb-saving reperfusion | 504  
    life-saving reperfusion | 504  
