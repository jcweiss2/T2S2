67 years old | 0
male | 0
admitted to the hospital | 0
left leg swelling | -168
cactus plant injury | -168
Primary Sclerosing Cholangitis | 0
mild Ulcerative Colitis | 0
deranged liver function tests | 0
presentation to ED | 0
left leg erythema | 0
left leg pain | 0
generally unwell | 0
paramedic assistance | 0
Blood Pressure 71/41mmHg | 0
Mean Arterial Pressure 48mmHg | 0
Respiratory Rate 36 breaths per minute | 0
Heart Rate 125 beats per minute | 0
sinus tachycardia | 0
Temperature 39°C | 0
Oxygen Saturation 86% | 0
admitted to ICU | 0
pH 7.15 | 0
PO2 84 | 0
HCO3 15 | 0
Lactate 7.6 | 0
Sodium 134 | 0
Urea 7.6 | 0
Creatinine 173 | 0
eGFR 27 | 0
White Cell Count 13.8 | 0
C-reactive protein 22 | 0
Hemoglobin 114 | 0
Platelet 81 | 0
Liver Function Test - Total Bilirubin 99 | 0
Alanine transaminase 61 | 0
Aspartate aminotransferase 83 | 0
Alkaline Phosphatase 96 | 0
Triple vasopressor support initiated | 0
Noradrenaline 20mcg/min | 0
Adrenaline 20mcg/min | 0
Vasopressin 0.04units/min | 0
Piperacillin-Tazobactam IV 4.5g | 0
Meropenem IV 2g | 0
Lincomycin IV 600mg | 0
Vancomycin IV 2g | 0
emergency left lower limb fasciotomy | 0
debridement | 0
below knee amputation | 0
necrotizing fasciitis | 0
LRINEC Score 5 | 0
extensive left foot and below knee tissue necrosis | 0
dishwasher fluid | 0
liquefied fat | 0
unviable skin and muscle | 0
histopathology | 0
post operatively | 24
transferred to ICU | 24
intubated | 24
possible re-exploration | 24
oliguria | 24
blood gas | 24
severe acidosis | 24
left internal jugular vascath insertion | 24
CRRT | 24
pH 7.28 | 24
Lactate 4.7 | 24
Sodium 130 | 24
Creatinine 206 | 24
Hemoglobin 89 | 24
Platelet 105 | 24
White Cell Count 17 | 24
C-reactive protein 78 | 24
International normalized ratio 2.2 | 24
Activated Partial Thromboplastin Time 150 | 24
Group B Streptococcus pneumoniae | 24
Ventilation sedation | 24
Propofol 170mg/hr | 24
Fentanyl 40mcg/hr | 24
CRRT on heparin circuit | 24
Renal dose 30ml/kg/hr | 24
Triple vasopressor support | 24
Noradrenaline 23mcg/min | 24
Adrenaline 18mcg/min | 24
Vasopressin 0.04units/min | 24
Antibiotics | 24
Meropenem IV 2g TDS | 24
Lincomycin IV 600mg TDS | 24
Vancomycin IV 2g BD | 24
Intravenous Immunoglobin G 100g | 24
taken back to theatre | 48
source control | 48
viability of the left stump | 48
no evidence of necrotic tissue | 48
Rapid Atrial Fibrillation | 48
HR 110bpm | 48
oliguric | 48
pH 7.40 | 48
Lactate 3.9 | 48
Sodium 131 | 48
Creatinine 116 | 48
White Cell Count 26 | 48
C-reactive protein 105 | 48
Procalcitonin 21.18 | 48
Hemoglobin 83 | 48
Platelet 63 | 48
INR 3.1 | 48
Fibrinogen 2.4 | 48
Echocardiography | 48
Moderate segmental left ventricular dysfunction | 48
Ejection Fraction 40-45% | 48
Dilated atria bilaterally | 48
Raised Right Atrial Pressure | 48
Amiodarone loading dose | 48
Amiodarone maintenance dose | 48
CRRT AN69 anti-inflammatory heparin laden adsorbing filter | 72
Citrate based anticoagulation circuit | 72
Sepsis Induced Coagulopathy | 72
bedside surgical debridement | 72
pH 7.31 | 72
Lactate 2.4 | 72
Sodium 135 | 72
Creatinine 79 | 72
White Cell Count 27 | 72
C-reactive protein 127 | 72
Hemoglobin 78 | 72
Platelet 50 | 72
INR 2.0 | 72
Histopathology | 72
NF | 72
Wound culture | 72
GBSPn | 72
Tissue culture | 72
GBSPn | 72
Vasopressor support weaning | 72
Noradrenaline 20mcg/min | 72
Adrenaline weaned off | 72
Vasopressin 2.4units/min | 72
oliguric | 96
Furosemide IV 250mg | 96
pH 7.36 | 96
Lactate 1.5 | 96
Sodium 130 | 96
Creatinine 116 | 96
White Cell Count 33 | 96
C-reactive protein 103 | 96
Procalcitonin 15.37 | 96
Hemoglobin 91 | 96
Platelet 53 | 96
INR 1.7 | 96
LFT - Bili 131 | 96
AST 127 | 96
ALP 121 | 96
Double inotropic support | 96
Noradrenaline 20mcg/min | 96
Vasopressin 2.4units/min | 96
fulminant hepatic failure | 120
encephalopathy | 120
refractory oliguria | 120
pH 7.39 | 120
Lactate 1.2 | 120
Sodium 134 | 120
Creatinine 124 | 120
White Cell Count 39.5 | 120
C-reactive protein 74 | 120
Hemoglobin 116 | 120
Platelet 49 | 120
INR 1.5 | 120
LFT- Bili 139 | 120
AST 69 | 120
ALT 97 | 120
ALP 140 | 120
Dual inotropic support | 120
Noradrenaline 20mcg/min | 120
Vasopressin weaned off | 120
ICU acquired weakness | 144
unarousable | 144
no response to noxious stimuli | 144
intubated | 144
ventilated | 144
Pressure Support Ventilation | 144
refractory oliguria | 144
pH 7.44 | 144
Lactate 1.1 | 144
White Cell Count 43.5 | 144
C-reactive protein 109 | 144
Hemoglobin 90 | 144
Platelet 57 | 144
INR 1.5 | 144
LFT - Bili 150 | 144
AST 95 | 144
ALP 154 | 144
Sedation weaned off | 144
Noradrenaline weaned off | 144
Antibiotic de-escalation | 144
Lincomycin ceased | 144
Vancomycin ceased | 144
Meropenem IV 2g TDS | 144
CRRT | 144
Hyper-Ammonium Therapy | 144
Rifaximin NGT 550mg BD | 144
Lactulose NGT 20ml TDS | 144
PRBCs transfusion | 144
jaundice | 168
Hypoactive delirium | 168
deeply sedated | 168
RASS -5 | 168
lateralizing signs | 168
CT Brain | 168
No acute intracranial pathology | 168
Ultrasound abdomen | 168
Acute Calculous Cholecystitis | 168
pH 7.44 | 168
Lactate 1.1 | 168
White Cell Count 44.3 | 168
C-reactive protein 109 | 168
Hemoglobin 129 | 168
Platelet 66 | 168
INR 1.3 | 168
LFT - Bili 235 | 168
AST 75 | 168
ALP 175 | 168
Conjugated Bilirubin 142 | 168
Meropenem IV 2g TDS | 168
CRRT | 168
Heparin circuit | 168
Anuria | 192
Hypotensive | 192
BP 71/33 | 192
MAP 51mmHg | 192
Febrile | 192
RAF | 192
HR 160 | 192
deterioration | 192
palliative care pathway | 192
deceased | 192
Troponin 616 | 192
Ammonia 158 | 192
LFT - Bili 352 | 192
AST 100 | 192
ALP 299 | 192
CRRT | 192
Renal recovery assessment | 192
Furosemide IV 250mg | 192
Acetazolamide IV 500mg | 192
Vasopressor support | 192
Noradrenaline 2.5mcg/min | 192
Lincomycin IV 600mg TDS | 192
Meropenem IV 2g TDS | 192
Digoxin IV 500mcg | 192
Metoprolol IV 15mg | 192