14 years old | 0
male | 0
near-drowning incident | -1
cardiopulmonary resuscitation (CPR) | -1
abdominal pain | 0
diffuse abrasions on his torso | 0
pneumoperitoneum | 0
pneumomediastinum | 0
intraabdominal free fluid | 0
hollow viscus perforation | 0
gross contamination with food debris | 1
total gastroesophageal junction (GEJ) disruption | 1
hemodynamically labile | 1
damage control procedure | 1
distal esophagus and the proximal stomach stapled closed | 1
discontinuity | 1
Four drains including a mediastinal drain and a gastrostomy (G) tube placed | 1
large bore nasogastric (NG) tube placed in the esophagus | 1
intraabdominal and mediastinal drains placed | 1
Fascia closed | 1
transferred to the Pediatric Intensive Care Unit (ICU) | 1
septic shock | 24
respiratory failure | 24
prolonged intubation | 24
deep venous thrombosis | 24
pulmonary embolism | 24
bilateral pleural effusions | 24
general deconditioning | 24
parenteral nutrition started | 24
extubated | 432
fluoroscopic evaluation demonstrated a leak in the esophagus | 432
stomach negative for leak | 432
enteral nutrition initiated via the G tube | 432
discharged | 1200
Ivor-Lewis distal esophagectomy with gastric pull-up for esophagogastric anastomosis | 2160
gastric conduit made along the lesser curvature | 2160
right thoracotomy performed | 2160
distal esophagus identified | 2160
tubularized portion of the stomach advanced into the chest | 2160
29 mm end-to-end anastomosis (EEA) stapler used to complete the esophagogastric anastomosis | 2160
leak test performed via upper endoscopy | 2160
jejunostomy tube placed | 2160
extubated | 2184
nutritionally supported with jejunostomy enteral feeds | 2184
esophagram showed no leak at the anastomosis | 2208
initiated on a liquid diet | 2208
discharged | 2220
tolerate a regular diet without difficulty | 2592
gaining weight and recovering well | 2592