39 years old | 0
male | 0
street vendor | 0
lives in Bangkok | 0
admitted to the hospital | 0
5-day fever | -120
myalgia | -120
breathlessness | -6
haemoptysis | -6
20-pack-year smoking | 0
high body temperature | 0
tachypnea | 0
respiratory distress | 0
no conjunctival suffusion | 0
no icteric sclera | 0
bilateral diffuse opacification pattern | 0
arterial blood gas | 0
pH 7.42 | 0
pCO2 35.7 | 0
pO2 55 | 0
SpO2 89% | 0
lactate 1.2 | 0
FiO2 1.0 | 0
normal complete blood count | 0
mild coagulopathy | 0
total bilirubin 1.51 | 0
alanine aminotransferase 48 | 0
creatinine 0.93 | 0
albumin 3.4 | 0
mild proteinuria | 0
microscopic haematuria | 0
Thai-Lepto score 8.5 | 0
intubation | 0
fresh blood suctioned | 0
admitted to intensive care unit | 0
APACHE II score 17 | 0
respiratory distress | 0
oxygen desaturation | 0
diffuse alveolar haemorrhage | 0
severe ARDS | 0
ventilator support | 0
lung-protective strategy | 0
sedations | 0
neuromuscular blockade | 0
cisatracurium | 0
propofol | 0
midazolam | 0
fentanyl | 0
ceftriaxone | 0
levofloxacin | 0
plasmapheresis | 2
intravenous pulse methylprednisolone | 2
VV-ECMO | 12
leptospirosis diagnosis | 24
leptospiral DNA detection | 24
anti-Leptospira IgM antibodies | 24
negative | 24
positive | 192
transthoracic echocardiography | 0
normal left ventricular size | 0
normal systolic function | 0
no vegetation | 0
haemoculture negative | 0
sputum culture negative | 0
anti-HIV negative | 0
anti-hepatitis C virus negative | 0
HBsAg negative | 0
anti-HBs negative | 0
anti-HBc negative | 0
Weil-Felix test negative | 0
OX 19 titre negative | 0
OX K titre negative | 0
OX 2 titre negative | 0
scrub typhus Ab negative | 0
murine typhus Ab negative | 0
dengue NS1 antigen negative | 0
dengue IgM negative | 0
dengue IgG positive | 0
influenza A/B/RSV rapid test negative | 0
RT-PCR negative | 0
respiratory virus 19 subtypes negative | 0
thin and thick blood films for malaria negative | 0
antinuclear antibodies negative | 0
CH50 44.9 | 0
C3 138 | 0
C4 53.4 | 0
renal function impaired | 0
returned to normal | 96
liver function test normal | 0
condition improved | 120
weaned off VV-ECMO | 120
withdrawal of VV-ECMO | 192
endotracheal tube | 192
discharged from intensive care unit | 240
discharged home | 336
follow-up | 8760
recovered | 8760