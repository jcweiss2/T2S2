26 years old | 0
female | 0
admitted to the hospital | 0
pregnant | 0
G1P1 | 0
no history of febrile urinary tract infection | 0
no history of flank pain | 0
no history of urolithiasis | 0
presented at 39 weeks of gestation | 0
normal vaginal delivery | 0
no complications | 0
prenatal care uneventful | 0
two screening urine analyses | -1680
two screening urine cultures | -1680
no evidence of infection | -1680
denied fever | 0
denied lower urinary tract symptoms | 0
sinus tachycardia | 0
maximal heart rate 142 beats per minute | 0
tachypnea | 0
dyspnea | 0
respiratory rate 20-24 breaths per minute | 0
hypotension | 0
maximal drop in systolic blood pressure 30 mmHg | 0
refractory to fluid boluses | 0
no fever | 0
normally contracted uterus | 0
no abnormalities noted in physical exam | 0
elevated white count 32,500/ml | 0
CT angiography of the chest | 0
suspected pulmonary embolism | 0
chest CT showed huge lesion occupying right kidney topography | 0
abdominal MRI | 0
pelvic MRI | 0
large multi-loculated multi-septated cystic mass | 0
mass arising from upper pole of right kidney | 0
mass measuring 19.0 × 15.5 × 16.5 cm | 0
mass abutting right hepatic lobe | 0
no definite infiltration | 0
mass effect on aorta | 0
mass effect on celiac axis | 0
mass effect on portal confluence | 0
mass effect on gallbladder | 0
mass effect on pancreas | 0
deviated to the left side | 0
no filling defect | 0
no obstructing stone | 0
differential diagnosis included multilocular cystic nephroma | 0
differential diagnosis included cystic renal carcinoma | 0
differential diagnosis included hydatid disease | 0
transferred to Intensive Care Unit | 0
broad-spectrum antibiotic coverage with meropenem | 0
broad-spectrum antibiotic coverage with vancomycin | 0
fever developed | 24
Tmax 39.1 °C | 24
slight worsening of hemodynamics | 24
lowest mean arterial pressure 59 mmHg | 24
decision to proceed with surgical exploration | 24
extended Chevron incision | 24
huge right kidney identified | 24
ascending colon medially retracted | 24
duodenum medially retracted | 24
perinephric tissue dissected anteriorly | 24
perinephric tissue dissected caudally | 24
extremely adherent posteriorly | 24
extremely adherent superomedially | 24
attempts to elevate kidney from psoas fascia | 24
eruption of large posterior cyst | 24
purulent foul-smelling grey-brown fluid spilled | 24
thorough irrigation of surgical field | 24
nephrectomy completed | 24
cleaning of surrounding suspicious-looking fat tissues | 24
postoperative period uneventful | 24
hemodynamics improved significantly after resection | 24
discharged 4 days postoperatively | 96
heart rate normalized | 96
blood pressure normalized | 96
afebrile at discharge | 96
urine culture grew multi-sensitive Escherichia coli | 96
pus culture grew multi-sensitive Escherichia coli | 96
gross specimen weight 1.26 kg | 96
kidney size 17 × 16 × 10 cm | 96
tan yellow mass | 96
soft mass | 96
cystic areas | 96
areas of necrosis | 96
histopathological examination revealed sheets of lipid-laden macrophages | 96
histopathological examination revealed histiocytes | 96
histopathological examination revealed multinucleated giant cells | 96
acute inflammation | 96
chronic inflammation | 96
involvement of renal parenchyma | 96
extension into perinephric fat | 96
extension into adrenal gland | 96
no evidence of hydatid cyst disease | 96
GMS stains negative for microorganisms | 96
PAS stains negative for microorganisms | 96
AFB stains negative for microorganisms | 96
xanthogranulomatous pyelonephritis | 96
seen 2 weeks after discharge | 336
vital signs within normal range | 336
wound clean | 336
no evidence of infection | 336
