43 years old | 0
female | 0
history of difficult-to-manage bronchial asthma | 0
hospitalized in the last 8 months on 10 occasions for acute exacerbations | -5736
hospitalized in the last 8 months on 10 occasions for asthmatic crisis | -5736
24-hour history of dry cough | -24
24-hour history of progressive dyspnea | -24
24-hour history of psychomotor agitation | -24
24-hour history of audible wheezing | -24
outpatient use of salbutamol | -24
outpatient use of ipratropium bromide | -24
admitted in critical condition | 0
diaphoretic | 0
tachycardic (heart rate 110 beats/minute) | 0
dyspneic with supraclavicular retractions | 0
respiratory rate of 30 breaths/minute | 0
ambient oxygen saturation 87% | 0
auscultation with abolished vesicular murmur in both lung fields | 0
Glasgow coma scale 12/15 | 0
arterial blood gases analysis revealed respiratory acidosis | 0
arterial blood gases analysis revealed hypoxemia | 0
pH: 7.21 | 0
PCO2: 66.5 | 0
PO2: 53.4 | 0
HCO3: 26.5 | 0
BE −2.8 | 0
SaO2 79.1% | 0
PaO2/FiO2: 178 | 0
invasive ventilatory support provided | 0
midazolam (loading dose 0.2 mg/kg) | 0
midazolam (maintenance dose 0.05 mg/kg/h) | 0
propofol (loading dose 1 mg/kg) | 0
propofol (maintenance dose 1 mg/kg/h) | 0
transferred to the ICU | 0
managed with hydrocortisone 100 mg IV every 8 hours | 0
managed with magnesium sulfate | 0
managed with antibiotics (piperacillin tazobactam and clarithromycin) | 0
infection as the cause of the asthmatic crisis | 0
day 2: short-term (48-hour) infusion of neuromuscular blocking agents (NMB) | 48
cisatracurium initial dose of 0.15 mg/kg | 48
cisatracurium maintenance dose of intermittent 0.03 mg/kg IV bolus | 48
train of 4 used to monitor paralysis maintaining a range of 1-2 | 48
day 4: improvement in ABG | 96
ventilatory weaning indicated | 96
suspending dual sedation | 96
suspending NMB | 96
light sedation with dexmedetomidine started | 96
day 6: GCS 15/15 | 144
weakness of the neck flexor muscles | 144
facial paresis | 144
could not move all 4 limbs | 144
muscular strength 1/5 in lower limbs | 144
muscular strength 2/5 in upper limbs | 144
flaccid hyporeflexia | 144
preserved sensitivity | 144
no alteration in cranial nerves | 144
assessed by neurology | 144
brain MRI requested | 144
cervical MRI requested | 144
study of cerebrospinal fluid requested | 144
brain MRI normal | 144
cervical MRI normal | 144
cerebrospinal fluid normal | 144
MRC score 37 points | 144
electromyography (EMG) performed | 144
EMG revealed signs of denervation | 144
EMG revealed signs of irritability (myopathic pattern) | 144
EMG revealed polyneuropathic compromise with axonal pattern in conduction velocity | 144
diagnosis of ICUAW confirmed | 144
physiotherapy started | 144
comprehensive rehabilitation started | 144
ventilator withdrawn achieved on day 10 | 240
hospital discharge | 720
30 days after admission | 720
MRC score of 55 points | 720
normal ABG control | 720
no acidosis | 720
no hypoxemia | 720
symptomatic resolution achieved | 720
