62 years old | 0
woman | 0
end-stage renal disease | -5760
regular haemodialysis via right-sided double-lumen tunnelled catheter | -5760
presented to emergency department | 0
progressive shortness of breath | -72
cough | -72
tachypneic | 0
temperature 37.7°C | 0
heart rate 110 beats per minute | 0
blood pressure 100/55 mmHg | 0
oxygen saturation 85% on room air | 0
clear lung fields | 0
pansystolic murmur over the right lower parasternal area | 0
computed tomography pulmonary angiography | 0
bilateral segmental and subsegmental pulmonary embolism | 0
polymerase chain reaction testing for SARS-CoV2 negative | 0
admitted to intensive care unit | 0
intravenous heparin infusion initiated | 0
hypotension | 48
blood pressure 70/40 mmHg | 48
transthoracic echocardiography | 48
dilated right side | 48
significant tricuspid regurgitation | 48
pulmonary artery systolic pressure 56 mmHg | 48
normal aortic valve | 48
ST-segment elevation in the inferolateral leads | 48
high-sensitive cardiac troponin-T increased | 48
coronary angiography | 48
total occlusion of the posterior descending artery | 48
multiple attempts for aspiration and balloon inflation failed | 48
relocated to ICU | 48
complete heart block | 72
temporary pacemaker insertion | 72
feverish | 72
temperature 38.9°C | 72
pus oozing from haemodialysis catheter site | 72
line sepsis diagnosed | 72
catheter removed | 72
blood culture revealed Methicillin-resistant Staphylococcus aureus | 72
catheter tip culture revealed Methicillin-resistant Staphylococcus aureus | 72
transesophageal echocardiography | 72
aortic valve vegetations | 72
acute severe aortic regurgitation | 72
right atrial appendage mass | 72
patent foramen ovale | 72
intravenous vancomycin initiated | 72
disturbed level of consciousness | 72
resistant shock | 72
mechanically ventilated | 72
intravenous inotropes increased | 72
extracorporeal membrane oxygenation system inserted | 72
died | 72
