29 years old | 0
primigravida | 0
32-week gestation | 0
admitted to the hospital | 0
sore throat | -240
high-grade fever | -240
abdominal pain | -240
cough | -240
progressive shortness of breath | -240
poor urine output | -48
decreased fetal movements | -48
uneventful pregnancy | -672
ultrasonography scan | -168
single live fetus | -168
normal biometry parameters | -168
tested for COVID-19 | -240
reverse transcriptase polymerase chain reaction assay | -240
COVID-19 suspect | 0
residence in containment zone | 0
investigated for COVID-19 | 0
RT-PCR assay | 0
negative COVID-19 test | 0
previous COVID-19 RT-PCR test | -240
negative previous COVID-19 test | -240
chest X-ray | 0
abdominal shielding | 0
minimal bilateral basal haziness | 0
prominent interstitial markings | 0
acute hypoxemic respiratory failure | 0
hypotension | 0
admitted to respiratory intensive care unit | 0
provisional diagnosis of community-acquired pneumonia | 0
septic shock | 0
inhaled oxygen supplementation | 0
intravenous fluids | 0
vasopressors | 0
broad-spectrum antibiotics | 0
fundal height corresponding to gestational age | 0
no fetal movements | 0
no fetal heart rate | 0
anemia | 0
leucocytosis | 0
mildly elevated C-reactive protein levels | 0
serum procalcitonin levels | 0
acute kidney injury | 0
mildly deranged liver function tests | 0
single intrauterine fetus | 0
no cardiac activity | 0
informed about intrauterine death | 0
high-risk consent for induction of labor | 0
delivery conducted | 24
stillborn male fetus | 24
no intrapartum adverse events | 24
no postpartum adverse events | 24
RT-PCR for COVID-19 negative | 0
Haemoglobin 11.2 | 0
Total leucocyte counts 20,300 | 0
Platelet counts 2.15 | 0
Serum Bilirubin 2.0 | 0
SGOT/SGPT 93/70 | 0
Serum Creatinine 2.5 | 0
C-Reactive Protein 9.8 | 0
S. Na+/K+ 132/4.3 | 0
Prothrombin Time 12.5 | 0
International Normalized Ratio 1.01 | 0
d-dimers 235 | 0
Blood culture sterile | 0
Urine culture sterile | 0
High vaginal swab culture sterile | 0
Work-up for Malaria negative | 0
Work-up for Dengue negative | 0
Work-up for Typhoid negative | 0
Work-up for Leptospira negative | 0
Work-up for H1N1 Influenza negative | 0
IgM Antibodies for Scrub typhus positive | 48
febrile illness | 0
work-up for tropical fevers | 48
peripheral smear negative | 48
antigen-based assays for malaria negative | 48
serology for dengue negative | 48
serology for leptospira negative | 48
serum Widal tests negative | 48
eschar detected | 48
doxycycline therapy started | 48
clinical response seen | 120
clinical–radiological parameters improved | 120
leukocyte counts normalized | 120
serum creatinine normalized | 120
vitals maintained without oxygen support | 168
discharged in stable condition | 168