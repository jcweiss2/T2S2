85 years old | 0
male | 0
admitted to the hospital | 0
melena | -3600
weakness | -3600
dizziness | -3600
abdominal aortic aneurysm repair | -2976
lower abdominal aorta-common iliac artery bifurcated stent implantation | -2976
gastrointestinal bleeding | -3360
tiredness | -2520
aspirin-induced mucosal injury | -2520
aspirin | -2520
blood transfusion | -2520
proton pump inhibitors | -2520
discharged | -2460
progressive fatigue | -1840
loss of appetite | -1840
weight loss | -1840
intermittent palpitation | -1840
intermittent fever | -1840
pneumonia | -1840
antibiotics | -1840
discharged | -1760
right back pain | -336
right knee movement restriction | -336
right leg swelling | -336
pale | 0
skinny | 0
body temperature | 0
pulse rate | 0
respiratory rate | 0
blood pressure | 0
abdomen soft | 0
nontender | 0
no palpable masses | 0
normal bowel sounds | 0
severe anemia | 0
white blood cell count | 0
granulocytes | 0
blood transfusion | 0
antibiotics | 0
computed tomography | 0
gas shadow | 0
thrombosis | 0
encapsulated fluid | 0
SAEF | 0
duodenoscopy | 0
fistula | 0
open surgery | 24
extraanatomic bypass | 24
infection | 24
intestinal erosion | 24
stent-induced infection | 24
excision of infected endograft | 24
aortic stent graft excision | 24
infrarenal abdominal aortic suture | 24
left common iliac artery ligation | 24
surgical debridement | 24
retroperitoneal abscess resolution | 24
drainage | 24
duodenal defect repair | 24
jejunal feeding tube placement | 24
operation time | 24
intensive care unit | 24
broad-spectrum intravenous antibiotics | 24
imipenem/cilastatin | 24
multiorgan function monitoring | 24
tissue from retroperitoneal abscess | 120
Enterococcus faecium | 120
Candida albicans | 120
vancomycin | 120
fluconazole | 120
hospital-acquired pneumonia | 240
bilateral pleural effusion | 240
heart failure | 240
wide-spectrum intravenous antibiotics | 240
cefoperazone/sulbactam | 240
fluid intake restriction | 240
progressive abdominal distension | 360
partial small-bowel obstruction | 360
postoperative intestinal adhesions | 360
fasting | 360
parenteral nutrition | 360
gastrointestinal decompression | 360
inhibition of gastric acid secretion | 360
oral paraffin fluid | 360
enema | 360
recovered | 720
discharged | 720