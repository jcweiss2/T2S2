Here is the extracted table of clinical events and timestamps:

COVID-19 pandemic | 0
respiratory system affected | 0
severe acute respiratory distress syndrome | 0
involvement of vital organs | 0
renal involvement | 0
acute kidney injury (AKI) | 0
pregnancy | 0
high-risk condition for COVID-19 disease | 0
deterioration | 0
secondary causes of AKI in pregnancy | 0
literature search | 0
PubMed search | 0
Scopus search | 0
Google Scholar search | 0
ScienceDirect search | 0
search strings used | 0
results retrieved | 0
studies screened | 0
studies short-listed | 0
studies excluded | 0
studies included | 0
AKI considered a surrogate marker of disease severity | 0
AKI predictor of outcome in terms of mortality | 0
AKI reported in 20%–40% of patients with COVID-19 | 0
intensive care | 0
RRT needed in 20% of affected patients | 0
incidence of AKI varies from 0.5% to 29% | 0
antenatal women high-risk group | 0
susceptibility to severe viral pneumonia increases | 0
changes in immune system | 0
pulmonary adaptations | 0
available literature undecided | 0
adverse maternal outcome in 3% of pregnant women | 0
associated comorbidities | 0
pregnancy leads to alterations in homeostatic mechanisms | 0
suppression of cellular immunity | 0
changes in hormonal milieu | 0
higher levels of progesterone and prostaglandins | 0
adverse outcome | 0
increased risk of spontaneous abortion | 0
hypertension | 0
prematurity | 0
adverse perinatal outcomes | 0
intrauterine death | 0
prognosis worst if disease acquired in last few weeks of gestation | 0
Asian or ethnic origin high-risk factor | 0
high body mass index high-risk factor | 0
mechanism of viral replication | 0
attachment of surface coronations to angiotensin-converting enzyme 2 receptors | 0
mitochondrial dysfunction | 0
acute tubular necrosis (ATN) | 0
protein reabsorption | 0
vacuole formation | 0
collapsing glomerulopathy | 0
protein exudates in Bowman's capsule | 0
etiology of renal damage multifactorial | 0
renal congestion secondary to right heart failure | 0
low cardiac output due to left ventricular dysfunction | 0
arterial hypotension | 0
renal damage due to direct tubular involvement | 0
cytokine storm caused by virus | 0
intravascular volume management essential | 0
fluid loss due to pyrexia and tachypnea | 0
positive fluid balance detrimental for lungs | 0
tremendous alteration in immune system | 0
immunosuppressed milieu during pregnancy | 0
exaggerated hormonal state | 0
increased predisposition to severe acute respiratory syndrome (SARS) infection | 0
subdued cellular immune response | 0
T helper cells (TH1 to TH2) shift | 0
altered hemodynamic state during pregnancy | 0
increased effect | 0
underlying kidney disease factor for deterioration | 0
development of complications | 0
mother and baby | 0
pregnant women had 51% increased risk of developing AKI | 0
independent of age and clinical comorbidities | 0
pregnancy increases risk of AKI | 0
case reports regarding AKI in pregnancy | 0
ATN in pregnancy with COVID-19 | 0
computed tomography of chest revealed ground-glass opacities | 0
consolidation in upper right lobe | 0
tachypnea | 0
rising creatinine levels | 0
respiratory and metabolic acidosis | 0
intubation | 0
dialytic support | 0
cesarean section | 0
dialysis 12 h before surgical intervention | 0
baby tested negative for COVID-19 | 0
oliguria | 0
diuretic use | 0
hemoperfusion | 0
resolution of ATN | 0
new-onset severe preeclampsia | 0
SARS-CoV-2-infected women | 0
termination of pregnancy | 0
preeclampsia as differential for acute liver injury | 0
placental histopathology | 0
vascular thrombi | 0
low-dose aspirin | 0
prevention of preeclampsia | 0
development of severe preeclampsia | 0
complicated by acute fatty liver of pregnancy (AFLP) | 0
hemolysis, elevated liver enzymes, and low platelets (HELLP) syndrome | 0
AKI | 0
endothelial injury | 0
common hallmark | 0
primary underlying pathogenetic mechanism | 0
COVID-19 infection | 0
endothelial disruption | 0
derangement in coagulation parameters | 0
thrombotic tendency | 0
preeclampsia | 0
worsening clinical picture | 0
renin-angiotensin-aldosterone system axis | 0
renal dysfunction | 0
recovery from COVID infection | 0
not affected by AKI | 0
similar picture in SARS CoV-induced AKI | 0
pregnancy-related renal and cardiovascular complications | 0
preeclampsia | 0
PR-AKI mostly occurs secondary to preeclampsia | 0
severe features | 0
HELLP | 0
other rare obstetric complications | 0
atypical hemolytic uremic syndrome | 0
thrombotic thrombocytopenic purpura | 0
AFLP | 0
outcome of CoV19 associated PR-AKI | 0
acute renal failure | 0
end-stage renal disease | 0
renal transplant | 0
maternal as well as perinatal outcome | 0
worse in women with PR-AKI | 0
prolonged ICU stay | 0
low birth weight | 0
stillbirth/perinatal death | 0
clinical features of preeclampsia and severe COVID-19 | 0
similar | 0
biochemical markers of preeclampsia | 0
fms-like tyrosine kinase-1 | 0
placental growth factor | 0
differentiate these two etiologies | 0
clinical manifestation of COVID-19-induced systemic inflammation | 0
similar to preeclampsia | 0
hallmark abnormal placentation | 0
resulting biochemical abnormalities | 0
lacking in COVID-19 infection | 0
prognosis guarded in women with PR-AKI | 0
coexisting COVID-19 sepsis | 0
management includes RRT | 0
ventilatory support | 0
optimal outcome | 0
clinical progression of AKI | 0
defined according to KDIGO criteria | 0
serum creatinine trends | 0
stage 1 AKI | 0
increase in serum creatinine by 0.3 mg/dl | 0
within 48 h | 0
or 1.5–1.9 times increase in serum creatinine | 0
from baseline | 0
within 7 days | 0
stage 2 AKI | 0
2.9 times increase in serum creatinine | 0
within 7 days | 0
stage 3 AKI | 0
3 times or more increase in serum creatinine | 0
within 7 days | 0
or initiation of RRT | 0
increased blood flow to kidneys in normal pregnancy | 0
changes in hormonal profile | 0
increase in plasma volume | 0
decreased net glomerular oncotic pressure | 0
slight physiological increase in renal size | 0
resulting changes in autoregulation | 0
increase in estimated glomerular filtration rate (eGFR) | 0
significantly | 0
peak of 40%–50% | 0
compared to nonpregnant levels | 0
lower serum creatinine | 0
urea | 0
uric acid levels | 0
cutoff for eGFR to diagnose AKI | 0
lower in pregnant individuals | 0
>0.8 mg/dL or >70.72 μmol/L | 0
data on COVID-19 | 0
severe AKI more frequently seen in affected patients | 0
respiratory failure | 0
AKI reported in 89.7% of patients | 0
required ventilatory support | 0
compared to 21.7% who did not | 0
65.5% of patients developed severe AKI | 0
stages 2 and 3 AKI | 0
compared with 6.7% of those who did not | 0
stage 1, 2, and 3 AKI developed | 0
in 46.5%, 22.4%, and 31.1% | 0
respectively | 0
83.6% stage 3 AKI | 0
reported in patients on mechanical ventilation | 0
almost all patients on ventilatory support required RRT | 0
median interval of 2 h | 0
from time of hospital admission | 0
about 20 min from mechanical ventilation | 0
to initiation of dialysis | 0
most patients underwent intermittent hemodialysis | 0
54% | 0
continuous RRT | 0
use of both modalities (RRT and intermittent hemodialysis) | 0
24.6% and 21.4% | 0
respectively | 0
mortality seen in 35% of those who developed AKI | 0
prognosis worse in those requiring RRT | 0
supportive care guidelines | 0
KDIGO | 0
avoidance of nephrotoxic agents | 0
serial estimation of serum creatinine | 0
monitoring of urine output | 0
early initiation of invasive hemodynamic monitoring | 0
critically ill patients | 0
prevention of occurrence | 0
reduction of severity of AKI | 0
prophylactic measures | 0
supportive ventilation | 0
avoidance of pulmonary damage | 0
high pressures | 0
hypervolemia | 0
right ventricle volume overload | 0
pulmonary edema | 0
renal congestion | 0
AKI | 0
clinical deterioration | 0
routine blood pressure checks | 0
all pregnant females affected with COVID-19 | 0
irrespective of prior history of elevated blood pressures | 0
predisposing factors for preeclampsia | 0
investigation of all pregnant females presenting with severe preeclampsia | 0
abnormal laboratory results | 0
COVID-19 test | 0
plain X-ray of chest | 0
obstetric complications | 0
affecting kidneys | 0
preeclampsia | 0
thrombotic microangiopathies | 0
acute cortical necrosis | 0
placental abruption | 0
puerperal sepsis | 0
acute pyelonephritis | 0
lupus flare in pregnancy | 0
systemic lupus erythematosus | 0
acute-on chronic kidney disease | 0
differential diagnoses | 0
SARS-CoV-2 sepsis | 0
associated renal dysfunction | 0
resulting pathology | 0
activation of renin-angiotensin-aldosterone pathway | 0
systemic manifestations | 0
hepatorenal failure | 0
platelet dysfunction | 0
coagulation disorders | 0
hypertension | 0
serial monitoring of arterial blood gases | 0
lactate levels | 0
markers of hypoxia induced renal | 0
liver as well as myocardial damage | 0
prophylactic measures | 0
preexisting mild renal dysfunction | 0
prevent further damage | 0
rising serum creatinine values | 0
delay or avoid progression to AKI | 0
advanced measures | 0
individualized cases | 0
clinical improvement not evident with supportive therapies | 0
evidence of immune dysregulation | 0
high levels of inflammatory cytokines | 0
high or medium cutoff membranes | 0
continuous venovenous hemodialysis | 0
clearance of damaging cytokines | 0
hemoperfusion | 0
sorbent cartridges | 0
beginning of cytokine storm | 0
prevention of cytokine-induced kidney damage | 0
intermittent RRT | 0
hyperkalemia | 0
metabolic acidosis | 0
KDIGO stage 3 | 0
pulmonary edema | 0
ARDS | 0
outcome measures | 0
urine output>500 ml/day | 0
normalization of other parameters | 0
CRRT | 0
do | 0
ECCO2R (RRT+) | 0
incorporates polypropylene membrane lung | 0
in series before filter in CRRT | 0
mechanical ventilation-dependent AKI | 0
VT returns to baseline | 0
pH>7.3 | 0
respiratory rate≤35/min | 0
ECMO | 0
oxygenator inserted in circuit of CVVH | 0
return line | 0
ARDS | 0
metabolic disorders | 0
fluid overload | 0
20% decrease of both creatinine and BUN | 0
effective UF volume of at least 35 mL/kg/h | 0
role of extracorporeal carbon dioxide removal (ECCO2R) | 0
hypercapnia | 0
respiratory acidosis | 0
AKI | 0
cases where escalation of ionotropic support is required | 0
sequential extracorporeal therapies | 0
removal of endotoxins and cytokines | 0
sepsis-like syndrome | 0
superadded bacterial infection | 0
beneficial | 0
hypovolemia | 0
diuretic agents | 0
avoidance | 0
especially in pregnancy | 0
intradialytic hypotension | 0
RRT | 0
fetal circulation | 0
renal-transplant recipients | 0
immunosuppressant drugs | 0
prevent graft rejection | 0
associated comorbidities | 0
predisposing to higher risk of severe COVID-19 infection | 0
outcome of COVID-19 in these patients | 0
usually favorable | 0
no cases reported in pregnancy after renal transplant | 0
modifications in immunosuppressive agents | 0
individualized | 0
according to disease severity | 0
level of immunosuppression | 0
required | 0
continuous monitoring of fetal parameters | 0
monitoring of drug levels | 0
renal parameters | 0
especially those with gastroenteritis | 0
resulting in diarrhea | 0
fluid depletion | 0
commonly seen in COVID-19 sepsis | 0
pregnancy a state of altered immunological response | 0
prevention of rejection of conceptus | 0
allow fetal development | 0
susceptible to various infections | 0
predisposing to various complications | 0
aggressively monitor these patients | 0
appropriate clinical examinations | 0
laboratory investigations | 0
low threshold for detection of various complications | 0
AKI associated with COVID-19 | 0
investigated in a timely manner | 0
literature search regarding AKI in COVID-19 in pregnancy | 0
performed on PubMed | 0
Scopus | 0
Google Scholar | 0
ScienceDirect | 0
relevant articles selected | 0
multiorgan failure secondary to SARS-CoV-2-induced cytokine storm | 0
similar to various important obstetrical complications | 0
preeclampsia | 0
placental abruption | 0
AFLP | 0
AKI secondary to other etiologies | 0
during pregnancy | 0
sepsis | 0
hemorrhage | 0
lupus flare | 0
COVID sepsis in this subset of pregnant women | 0
urgent supportive care | 0
evaluation for inflammatory markers | 0
imaging | 0
differentiation of covid infection from other obstetrical conditions | 0
termination of pregnancy | 0
good maternal and neonatal outcome | 0