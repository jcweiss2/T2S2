58 years old | 0
female | 0
altered mental status | 0
difficulty breathing | 0
intermittent weakness | -720
fever | -720
rash | -720
tick exposures | -720
hypotensive | 0
hypoxic | 0
intubated | 0
vasopressors initiated | 0
creatinine of 203.32 μmol/L | 0
albumin of 17 g/L | 0
aspartate aminotransferase of 110 unit/L | 0
white blood cell count of 3.4 × 10^9/L | 0
hemoglobin level of 80 g/L | 0
hematocrit level of 26% | 0
platelet count of 36 × 10^9/L | 0
admitted to the intensive care unit | 0
lumbar puncture performed | 0
urinalysis sent | 0
urine culture sent | 0
blood culture sent | 0
blood test for tick-borne infections sent | 0
treated for septic shock with acute respiratory distress syndrome | 0
vancomycin administered | 0
cefepime administered | 0
doxycycline administered | 0
chest x-ray showed bilateral diffuse infiltrates | 0
acute respiratory distress syndrome management protocol started | 0
troponin level checked | 0
troponin level of 10 ng/mL | 0
electrocardiogram (ECG) performed | 0
transthoracic echocardiogram performed | 0
left ventricular ejection fraction (LVEF) of 55% to 60% | 0
left ventricular end-systolic volume index of 26 mL/m2 | 0
left ventricular end-diastolic volume index 67 mL/m2 | 0
normal wall motion | 0
elevated troponin thought to be a type 2 myocardial infarction | 0
troponin I level increased to > 40 ng/mL | 24
telemetry showed episodes of nonsustained ventricular tachycardia (NSVT) | 24
repeat ECG revealed low-voltage QRS with ST-segment elevation | 24
coronary angiography showed normal coronary arteries | 24
blood and urine cultures remained negative for 5 days | 120
urinalysis was unremarkable except for elevated myoglobin levels | 120
polymerase chain reaction (PCR) was negative for herpes simplex virus and cytomegalovirus | 120
Ehrlichia chaffeensis PCR from her blood sample was positive | 120
hepatitis panel showed no immunity or prior exposure to hepatitis A, B, or C | 120
Rocky Mountain Spotted Fever titers showed elevated levels of immunoglobulin-G antibody (Ab) | 120
vancomycin and cefepime stopped | 120
doxycycline continued | 120
respiratory status improved | 192
extubated | 192
frequent premature ventricular contractions | 192
multiple episodes of NSVT | 192
high suspicion for myocarditis | 192
cardiac magnetic resonance imaging performed | 192
global hypokinesis | 192
LVEF of 32% | 192
left ventricular mass of 45 g/m2 | 192
delayed enhancement in multiple areas of the myocardium and pericardium consistent with myopericarditis | 192
carvedilol administered | 192
lisinopril administered | 192
discharged to inpatient rehabilitation | 384
cardiomyopathy persisted | 4320
repeat transthoracic echocardiogram revealed an LVEF of 25% | 4320
repeat ECG revealed an improvement in QRS voltages | 4320
intermittent episodes of NSVT | 4320
amiodarone administered | 4320
cardioverter-defibrillator implanted | 4320
admissions for acute heart failure exacerbation | 8760