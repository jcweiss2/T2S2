61 years old | 0
Indigenous | 0
man | 0
presented to our hospital | 0
fever | -96
malaise | -96
cough | -96
breathlessness | -96
seropositive rheumatoid arthritis | -96
cutaneous lupus erythematosus | -96
emphysema | -96
ischaemic heart disease | -96
functional hyposplenism | -96
weekly subcutaneous etanercept | -12960
methotrexate | -12960
hydroxychloroquine | -12960
anemia | -1440
allergy to sulfanilamide | -87600
blistering skin rash | -87600
cigarette smoker | 0
not consumed alcohol | -26280
never injected intravenous drugs | 0
no history of recent gardening | 0
no history of soil exposure | 0
heart rate 104 beats per minute | 0
respiratory rate 24 breaths per minute | 0
blood pressure 101/56 mmHg | 0
oxygen saturation 97% | 0
temperature 39.7 °C | 0
hypopigmented rash | 0
right upper chest bronchial breath sounds | 0
crepitations | 0
mild left flank tenderness | 0
normocytic anemia | 0
leucocytosis | 0
neutrophilia | 0
acute kidney injury | 0
plain chest radiograph | 0
right upper lobe opacification | 0
left heart border opacification | 0
community-acquired pneumonia | 0
intravenous ceftriaxone | 0
intravenous gentamicin | 0
oral doxycycline | 0
deteriorated | 0
hypoxia | 0
hypotension | 0
hyperlactatemia | 0
oxygen via high-flow nasal-prongs | 0
intravenous noradrenaline | 0
intravenous meropenem | 0
intravenous vancomycin | 0
oral azithromycin | 0
transferred to the intensive care unit | 0
chest computerized tomography | 0
pulmonary infiltrates | 0
pneumonia | 0
no definite features of abscess formation | 0
no definite features of empyema | 0
no definite features of cavitation | 0
blood cultures collected at presentation | 0
Gram-negative bacilli | 0
Acinetobacter baumannii complex | 0
sensitive to meropenem | 0
sensitive to ceftazidime | 0
sensitive to co-trimoxazole | 0
sensitive to gentamicin | 0
second set of blood cultures | 72
Burkholderia pseudomallei | 72
sensitive to meropenem | 72
sensitive to co-trimoxazole | 72
sensitive to doxycycline | 72
isolates re-assessed for error | 72
no errors identified | 72
blood group testing | 72
sputum samples unable to be collected | 72
improved clinically | 168
discharged from ICU | 168
no ongoing oxygen requirement | 168
subsequent blood cultures | 168
no growth | 168
intravenous ceftazidime | 168
diagnosis of melioidosis | 168
CT scan of abdomen and pelvis | 168
visceral disease excluded | 168
L3/L4 discitis | 168
vertebral osteomyelitis | 168
lumbar spine magnetic resonance imaging | 168
peripherally inserted central catheter | 168
intravenous ceftazidime via elastomeric infusion | 168
etanercept withheld | 168
inflammatory arthritis managed | 168
simple analgesia | 168
low-dose corticosteroids | 168
concurrent oral TMP/SMX | 168
initially well tolerated | 168
oral TMP/SMX | 168
fixed drug eruption | 504
cessation of TMP/SMX | 504
change to doxycycline | 504
hyperlactatemia |0
oxygen via high-flow nasal-prongs |0
intravenous noradrenaline |0
intravenous meropenem |0
intravenous vancomycin |0
oral azithromycin |0
transferred to the intensive care unit |0
chest computerized tomography |0
pulmonary infiltrates |0
pneumonia |0
no definite features of abscess formation |0
no definite features of empyema |0
no definite features of cavitation |0
blood cultures collected at presentation |0
Gram-negative bacilli |0
Acinetobacter baumannii complex |0
sensitive to meropenem |0
sensitive to ceftazidime |0
sensitive to co-trimoxazole |0
sensitive to gentamicin |0
second set of blood cultures |72
Burkholderia pseudomallei |72
sensitive to meropenem |72
sensitive to co-trimoxazole |72
sensitive to doxycycline |72
isolates re-assessed for error |72
no errors identified |72
blood group testing |72
sputum samples unable to be collected |72
improved clinically |168
discharged from ICU |168
no ongoing oxygen requirement |168
subsequent blood cultures |168
no growth |168
intravenous ceftazidime |168
diagnosis of melioidosis |168
CT scan of abdomen and pelvis |168
visceral disease excluded |168
L3/L4 discitis |168
vertebral osteomyelitis |168
lumbar spine magnetic resonance imaging |168
peripherally inserted central catheter |168
intravenous ceftazidime via elastomeric infusion |168
etanercept withheld |168
inflammatory arthritis managed |168
simple analgesia |168
low-dose corticosteroids |168
concurrent oral TMP/SMX |168
initially well tolerated |168
oral TMP/SMX |168
fixed drug eruption |504
cessation of TMP/SMX |504
change to doxycycline |504
