64 years old | 0
    woman | 0
    poorly controlled diabetes mellitus | 0
    relapsing urinary tract infection | 0
    admitted to the intensive care unit | 0
    lower back pain | 0
    acute respiratory failure | 0
    septic shock | 0
    travelled to India | -1440
    nonsteroidal anti-inflammatory drugs | -1440
    no evidence for pneumonia | 0
    no ARDS | 0
    initial echocardiography | 0
    severe acute cor pulmonale | 0
    akinesia of the interventricular septum | 0
    electrocardiogram | 0
    transient ST segment elevation in the anteroseptal leads | 0
    coronary angiogram | 0
    atheromatous coronary arteries | 0
    no severe stenosis | 0
    abdominal computed tomography | 0
    gas collection in the parenchyma | 0
    gas collection in the perinephric space | 0
    gas in vein of the left kidney | 0
    control echocardiography at day-1 | 24
    no more acute cor pulmonale | 24
    no akinesia | 24
    emphysematous pyelonephritis | 0
    complicated by septic shock | 0
    multiple gas emboli in the pulmonary artery | 0
    transient cor pulmonale | 0
    gas emboli in the coronary artery | 0
    transient acute coronary syndrome | 0
    Klebsiella pneumoniae isolated in blood | 0
    Klebsiella pneumoniae isolated in urine | 0
    Klebsiella pneumoniae isolated in kidney cultures | 0
    treated with antimicrobials | 0
    treated with nephrectomy | 0
    favorable course | 0