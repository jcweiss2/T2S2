male | 0 | 0 
25-year-old mother | 0 | 0 
primigravida | 0 | 0 
uncomplicated pregnancy | -280 | 0 
spontaneous onset of labor | -1 | 0 
fetal distress | -1 | 0 
ventouse-assisted delivery | 0 | 0 
birth weight 3940 grams | 0 | 0 
resuscitation with mask ventilation | 0 | 0 
intubated | 0.13 | 0.13 
transferred to NICU | 0.13 | 0.13 
synchronized intermittent positive pressure ventilation (SIPPV) | 0.13 | 13.5 
gentamicin 4 mg/kg 24-hourly | 0 | 120 
benzyl penicillin 60 mg/kg 12-hourly | 0 | 13.5 
neutropenia | 18 | 18 
elevated inflammatory markers | 18 | 18 
C-reactive protein (CRP; 60 mg/L) | 18 | 18 
procalcitonin (68.55 µg/L) | 18 | 18 
lumbar puncture | 23 | 23 
normal cell count | 23 | 23 
negative for pathogens | 23 | 23 
placental surface eSwab | 23 | 23 
Gram-negative diplococci | 23 | 23 
Neisseria meningitidis | 23 | 23 
molecular testing | 23 | 23 
real-time PCR assay | 23 | 23 
N. meningitidis genogroup W DNA | 5.5 | 5.5 
blood cultures negative | 0.48 | 0.48 
benzylpenicillin dosage decreased | 13.5 | 13.5 
cefotaxime 50 mg/kg 12-hourly | 13.5 | 120 
elevated leucocyte count | -2.5 | -2.5 
neutrophil count of 18.1×10^9/L | -2.5 | -2.5 
maternal well after birth | 0 | 192 
baby improved | 13.5 | 192 
discharged home | 192 | 192 
contact tracing | 192 | 192 
chemoprophylaxis with ciprofloxacin | 192 | 192 
quadrivalent conjugate meningococcal vaccine | 192 | 192 
funisitis | -1 | 0 
chorioamnionitis | -1 | 0 
materno-fetal transmission | -1 | 0 
early-onset neonatal sepsis | 0 | 192 
invasive meningococcal disease (IMD) | 0 | 192 
N. meningitidis W CC11 | 0 | 192 
urethritis | -10080 | -10080 
Australia IMD rates due to N. meningitidis W | -10080 | 0 
case fatality rates | -10080 | 0 
public health concern | 192 | 192 
treatment and control measures | 192 | 192 
written consent | 0 | 0 
financial support | 0 | 0 
potential conflicts of interest | 0 | 0 
author contributions | 0 | 0 
laboratory and clinical work | 0 | 192 
diagnostic testing | 0 | 192 
clinical management | 0 | 192 
manuscript writing | 0 | 192 
oversight of the project | 0 | 192