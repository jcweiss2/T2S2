38 years old | 0
woman | 0
gravida 2 para 1 | 0
presented acutely at 9+0 weeks of gestation | 0
heavy vaginal bleeding | 0
signs consistent with hypovolaemic shock | 0
obstetric history included one caesarean section for breech presentation three years earlier | -8760
serial ultrasounds between 5 and 8 weeks of gestation | -4320
viable intrauterine pregnancy | 0
concurrent cystic structure in the lower uterine cavity at the site of the caesarean scar | 0
clinical concern for a heterotopic pregnancy with rupture of the non-viable caesarean scar pregnancy | 0
patient remained unstable despite resuscitation | 0
emergency examination under anaesthesia | 0
dilation and curettage | 0
laparotomy | 0
hysterectomy | 0
expressed a strong desire to preserve the viable intrauterine pregnancy and her uterus | 0
repeat bedside ultrasound showed a viable fundal intrauterine pregnancy | 0
lower uterine segment distension | 0
large blood clot | 0
ongoing bleeding | 0
ultrasound-guided suction curettage of the lower segment | 0
removal of thrombus and products of conception | 0
Foley catheter inserted into the uterus | 0
Foley catheter inflated to 70 ml | 0
Foley catheter placed under traction | 0
persistent bleeding | 0
decision to proceed with a laparotomy | 0
intra-operatively no evidence of uterine scar rupture | 0
bilateral uterine artery ligation performed | 0
significant reduction in vaginal bleeding | 0
massive transfusion intra-operatively with six units packed red blood cells | 0
four units of fresh frozen plasma | 0
haemoglobin 96 g/L at the close of the case | 0
admitted to the intensive care unit | 0
Foley catheter removed on day 3 post-operatively | 72
ultrasound at 9+4 weeks of gestation | 96
single live fetus | 96
heterogenous area in the lower segment of the uterus measuring 61×46×45 mm | 96
anterior myometrium intact throughout its length | 96
no free fluid in the pouch of Douglas | 96
discharged home on day 6 post-operatively | 144
serial ultrasounds between 11 and 20 weeks of gestation | 240
gradual resolution of the clot at the lower uterine segment to 14x11x5mm | 240
at 27+0 weeks of gestation | 4536
shortened cervix to 20 mm | 4536
commenced on vaginal progesterone | 4536
serial ultrasound at 27+6 weeks of gestation | 4608
cervical shortening to 11 mm | 4608
preterm rupture of membranes | 4608
emergency lower-segment caesarean section at 28+1 weeks of gestation | 4800
complete course of antenatal steroids | 4800
magnesium sulphate | 4800
caesarean section uncomplicated | 4800
liveborn male infant (1200 g, 56% for gestation) | 4800
admitted to the neonatal intensive care unit | 4800
neonate died on day 3 of life | 4824
extreme prematurity | 4824
respiratory distress syndrome | 4824
bilateral grade three intraventricular haemorrhages | 4824
two years later | 17520
spontaneously conceived pregnancy | 17520
complicated by placenta percreta | 17520
elective laparotomy | 17520
classical caesarean section | 17520
total abdominal hysterectomy at 34 weeks of gestation | 17520
complicated by a 6000 ml intra-operative haemorrhage | 17520
neonate born in good condition | 17520
admitted to the neonatal high-dependency unit for respiratory support | 17520
admitted to the intensive care unit for supportive care | 17520
discharged home in a good condition on day 11 post-operatively | 17520
