55 years old | 0
male | 0
admitted to the hospital | 0
severe watery diarrhoea | -576
opening his bowels 8–9 times in 24 h | -576
no other significant symptoms | -576
normal colonoscopy | -72
no past medical or surgical history | 0
no regular medications | 0
no significant family history | 0
non-smoker | 0
lethargic | 0
clinically dehydrated | 0
eGFR of 14 mL/min/1.73 m2 | 0
creatinine of 381 μmol/L | 0
serum potassium low at 2.5 mmol/L | 0
serum calcium elevated at 2.88 mmol/L | 0
normal anion gap metabolic acidosis | 0
pH of 7.16 | 0
base excess of −14.2 mmol/L | 0
normal lactate at 0.8 mmol/L | 0
inflammatory markers within the normal range | 0
coeliac serology negative | 0
vasculitis screen negative | 0
stool cultures negative | 0
admitted to the intensive care unit | 0
central potassium replacement | 0
aggressive rehydration with i.v. fluids | 0
parenteral nutrition commenced | 0
contrast-enhanced CT scan of the abdomen | 24
32-mm heterogenous mass in the pancreatic body | 24
multiple hypo-attenuating lesions throughout the liver parenchyma | 24
liver metastases | 24
radiological stage T2 N0 M1 | 24
fasting serum gut hormone profile sent | 24
somatostatin level 116 pmol/L | 24
gastrin level 47 pmol/L | 24
glucagon level 66 pmol/L | 24
chromogranin A level 223 pmol/L | 24
C terminal end chromogranin B level >4500 pmol/L | 24
VIP level 211 pmol/L | 24
PP level 6928 pmol/L | 24
ultrasound-guided core biopsy of a segment V liver lesion | 48
histology reported as mainly necrotic tissue | 48
viable tumour cells expressed epithelial marker CK8/18 | 48
viable tumour cells expressed neuroendocrine markers synaptophysin and CD56 | 48
chromogranin A expression negative | 48
Ki-67 proliferation index 2.9% | 48
p53 WT expression | 48
i.v. somatostatin analogue infusion initiated | 48
octreotide infusion at 12.5 µg/h | 48
diarrhoea settled completely | 48
renal function failed to improve | 72
spiking high temperatures | 72
inflammatory markers increased | 72
repeat CT showed significant amounts of intra-intestinal fluid | 72
blood cultures positive for K lebsiella and Enterococcus | 72
autonecrosis of the pancreatic primary and liver lesions | 72
treated for bowel bacteria overgrowth sepsis | 72
ultrafiltration commenced | 96
renal function improved significantly | 120
inflammatory markers settled | 120
stepped down to the ward | 120
discharged | 720
eGFR at discharge 54 mL/min/1.73 m2 | 720
Gallium-68 DOTA-TATE PET CT | 720
MRI of liver | 720
stable disease | 720
good response to SSA | 720
no evidence of disease beyond pancreas and liver | 720
lanreotide injections | 720
plan to proceed to surgical resection of primary tumour | 720
plan to debulk liver lesions | 720