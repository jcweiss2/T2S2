48 years old|0
Caucasian|0
female|0
found unresponsive at the scene of a house fire|0
burns to the face|0
<1% total body surface area (BSA)|0
inhalation injury|0
intubated via endotracheal tube|-0
transferred to our burn center|0
initial bronchoscopy showed diffuse carbonaceous sputum|-0
pale friable mucosa extending throughout the airways|-0
intubated for airway protection|0
required adequate sedation|0
neuromuscular blockade|0
diagnosis of severe depression with psychotic features|0
home medications included paliperidone palmitate 234 mg once monthly|0
paliperidone 6 mg by mouth daily|0
citalopram 40 mg by mouth daily|0
trazodone 150 mg by mouth at bedtime|0
risperidone 2 mg by mouth twice daily|0
clonazepam 1 mg by mouth twice daily|0
no known drug allergies|0
chronic smoker|0
substance abuser|0
urine drug screen was negative|0
mild leukocytosis|0
white blood cell count 15.8 k/mm3|0
afebrile|0
normotensive|0
adequate urine output (>0.5 mL/kg/hr)|0
evidence of acute respiratory distress syndrome (ARDS)|0
ratio of partial pressure arterial oxygen and fraction of inspired oxygen of less than 200|0
started on pressure control ventilation|0
tracheostomy was performed on the second hospital day (HD)|48
post-operatively became febrile|48
associated tachycardia|48
HD 5 expressed thick yellow secretions during suctioning|120
diffuse rhonchi|120
worsening right-sided, patchy infiltrate seen on chest X-ray|120
BAL culture on HD 6 revealed gram-positive cocci in clusters|144
blood cultures obtained on HD 4 grew Gram-positive cocci in clusters|96
started on empiric vancomycin and cefepime on HD 6|144
aggressive vancomycin dosing schedule (1750 mg IV every 6 h)|144
adequate, supratherapeutic, vancomycin trough concentrations of 26 mg/L|144
clinical status did not improve|144
continued febrile|144
tachycardic|144
increased ventilatory support|144
increased oxygenation requirements|144
repeat urine cultures on HD 5 were negative|120
repeat blood cultures on HD 5 were negative|120
Gram-positive pathogen identified as MRSA|120
repeat bronchoscopy on HD 10 demonstrated mild improvement in secretions|240
Gram-stain from the BAL yielded growth in culture of >110,000 CFU/mL MRSA|240
vancomycin MIC of 2 mg/L|240
deteriorating clinical status on HD 10|240
decision to modify antibiotic regimen|240
MRSA bacteremia and/or pneumonia|240
vancomycin MIC of ≥2 mg/L|240
linezolid not employed due to drug-drug interactions|240
initiate ceftaroline fosamil|240
ceftaroline MIC of 0.5 mg/L|240
ceftaroline regimen 600 mg IV every 8 h|240
became afebrile 48 h after initiation of ceftaroline|240
remained afebrile for the length of the hospital stay|240
rapid clinical improvement|240
weaned from the ventilator on HD 22|528
decannulated 2 days later|576
psychiatric illness|0
auditory/visual hallucinations|0
hospital discharge delayed|1152
serum concentrations of ceftaroline obtained for PK characterization|240
ceftaroline levels 30 min post-infusion: 21.9 mg/L|240
ceftaroline levels 2 h later: 7.3 mg/L|240
ceftaroline levels 30 min prior to next dose: 4.2 mg/L|240
ceftaroline half-life 1.5 h|240
ceftaroline Cmax 27.5 mg/L|240
ceftaroline Cmin 1.69 mg/L|240
ceftaroline Vd 0.42 L/kg|240
ceftaroline AUC0–τ 87.6 µg h/mL|240
ceftaroline T > MIC 8 h|240
ceftaroline clearance 10 L/h|240
continued for total of 14 days|240
completed ceftaroline therapy|240
resolved signs and symptoms of infection|240
no reported toxicity from antimicrobial therapy|240
liberated from mechanical ventilation|576
discharged on HD 48|1152
