65 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
admitted to the hospital | 0 | 0 | Factual
abdominal pain | -2160 | 0 | Factual
pancreatic head lesion | -2160 | 0 | Factual
history of stage IIIA lung cancer | -6480 | -6480 | Factual
smoking history | -6480 | 0 | Factual
hypertension | -6480 | 0 | Factual
hypothyroidism | -6480 | 0 | Factual
dyslipidemia | -6480 | 0 | Factual
spiculated suprahilar RUL nodule | -6480 | -6480 | Factual
lung-RADS 4X | -6480 | -6480 | Factual
PET/CT scan | -6480 | -6480 | Factual
bronchoscopy-attained tissue sample | -6480 | -6480 | Factual
NSCLC | -6480 | -6480 | Factual
adenocarcinoma | -6480 | -6480 | Factual
lymph node sampling | -6480 | -6480 | Factual
stage IIIA lung adenocarcinoma | -6480 | -6480 | Factual
program death ligand-1 expression | -6480 | -6480 | Factual
surgical resection | -6480 | -6480 | Negated
carboplatin | -5040 | -4320 | Factual
paclitaxel | -5040 | -4320 | Factual
radiation therapy | -5040 | -4320 | Factual
CT scan | -4320 | -4320 | Factual
decrease in RUL mass | -4320 | -4320 | Factual
adjuvant immunotherapy | -3960 | -3744 | Factual
durvalumab | -3960 | -3744 | Factual
pneumonitis | -3744 | -3744 | Factual
steroid taper | -3744 | -3744 | Factual
staging chest CT | -3744 | -3744 | Factual
increase in RUL mass | -3744 | -3744 | Factual
follow-up chest CT | -2160 | -2160 | Factual
increase in RUL mass | -2160 | -2160 | Factual
thoracic, abdominal, and pelvic CT scan | -1440 | -1440 | Factual
no distant metastasis | -1440 | -1440 | Factual
stable lung nodules | -1440 | -1440 | Factual
chest CT scans | -720 | -720 | Factual
stable appearance of lung nodules | -720 | -720 | Factual
post-radiation changes | -720 | -720 | Factual
epigastric pain | -120 | 0 | Factual
constipation | -120 | 0 | Factual
loss of appetite | -120 | 0 | Factual
weight loss | -120 | 0 | Factual
abdominal and pelvic CT scan | 0 | 0 | Factual
pancreatic head mass | 0 | 0 | Factual
pancreatic ductal dilatation | 0 | 0 | Factual
gastroenterology referral | 0 | 0 | Factual
endoscopic ultra-sound-guided biopsy | 24 | 24 | Factual
tumor cells | 24 | 24 | Factual
nuclear pleomorphism | 24 | 24 | Factual
prominent nucleoli | 24 | 24 | Factual
irregular nuclear contours | 24 | 24 | Factual
coarse chromatin | 24 | 24 | Factual
CK7 | 24 | 24 | Factual
TTF-1 | 24 | 24 | Factual
Napsin-A | 24 | 24 | Factual
CDX-2 | 24 | 24 | Negated
KOC | 24 | 24 | Negated
synaptophysin | 24 | 24 | Negated
Smad-4 | 24 | 24 | Factual
lung adenocarcinoma | 24 | 24 | Factual
AST | 24 | 24 | Factual
ALT | 24 | 24 | Factual
ALP | 24 | 24 | Factual
total bilirubin | 24 | 24 | Factual
direct bilirubin | 24 | 24 | Factual
CA 19.9 | 24 | 24 | Factual
PET/CT scan | 168 | 168 | Factual
fluorodeoxyglucose-avid mass | 168 | 168 | Factual
SUV max | 168 | 168 | Factual
brain MRI scan | 168 | 168 | Factual
no intracranial metastasis | 168 | 168 | Factual
palliative radiation therapy | 336 | 336 | Factual
carboplatin | 336 | 336 | Factual
pemetrexed | 336 | 336 | Factual
combination chemotherapy | 336 | 336 | Factual
generalized weakness | 720 | 720 | Factual
dyspnea | 720 | 720 | Factual
electrolyte derangements | 720 | 720 | Factual
acute anemia | 720 | 720 | Factual
hemoglobin nadir | 720 | 720 | Factual
transfusion | 720 | 720 | Factual
CT scan of the chest | 720 | 720 | Factual
new left lower lobe nodule | 720 | 720 | Factual
staging PET/CT scan | 1008 | 1008 | Factual
decreased metabolic activity | 1008 | 1008 | Factual
metabolic activity | 1008 | 1008 | Factual
fatigue | 1008 | 1008 | Factual
treatment discontinuation | 1008 | 1008 | Factual
pulmonology clinic | 1176 | 1176 | Factual
rapid response | 1176 | 1176 | Factual
oxygen saturation | 1176 | 1176 | Factual
accessory muscles | 1176 | 1176 | Factual
blood pressure | 1176 | 1176 | Factual
heart rate | 1176 | 1176 | Factual
increased dyspnea | 1176 | 1176 | Factual
cough | 1176 | 1176 | Factual
generalized weakness | 1176 | 1176 | Factual
emergency department | 1176 | 1176 | Factual
hospital admission | 1176 | 1176 | Factual
imaging studies | 1176 | 1176 | Factual
right lung consolidation | 1176 | 1176 | Factual
loculated pleural effusion | 1176 | 1176 | Factual
acute hypoxic respiratory failure | 1176 | 1176 | Factual
sepsis | 1176 | 1176 | Factual
pneumonia | 1176 | 1176 | Factual
broad-spectrum antibiotics | 1176 | 1176 | Factual
vancomycin | 1176 | 1176 | Factual
azithromycin | 1176 | 1176 | Factual
cefepime | 1176 | 1176 | Factual
oxygen supplementation | 1176 | 1176 | Factual
bilevel-positive airway pressure | 1176 | 1176 | Factual
altered mentation | 1248 | 1248 | Factual
worsening hypoxemia | 1248 | 1248 | Factual
vasopressor support | 1248 | 1248 | Factual
palliative medicine team | 1248 | 1248 | Factual
inpatient hospice care | 1248 | 1248 | Factual
death | 1260 | 1260 | Factual