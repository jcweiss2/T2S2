70 years old | 0
male | 0
farmer | 0
presented to the emergency department | 0
high-grade fever | -120
generalized body ache | -120
headache | -120
altered sensorium | -24
joint pains | 0
epigastric pain | 0
no other comorbidities | 0
no history of drug addiction | 0
no history of intoxication | 0
inguinal lymphadenopathy | 0
mild generalized rash | 0
no eschar | 0
hemodynamically stable | 0
disoriented | 0
no focal neurological deficit | 0
no neck rigidity | 0
acute febrile illness | 0
undifferentiated fever | 0
negative for malaria | 0
negative for dengue | 0
negative for typhoid | 0
negative for leptospira | 0
scrub typhus antigen card positive | 0
scrub IgM positive | 0
scrub typhus | 0
sterile blood cultures | 0
sterile other body fluid cultures | 0
leukocytosis (15,800/cc) | 0
mild hyperbilirubinemia | 0
transaminitis | 0
total bilirubin 3.6 mg/dL | 0
direct bilirubin 2.6 mg/dL | 0
serum glutamic oxaloacetic transaminase 116 U/L | 0
serum glutamic pyruvic transaminase 178 U/L | 0
slightly raised international normalized ratio (1.56) | 0
negative viral markers for hepatitis B antigen | 0
negative viral markers for hepatitis C antibody | 0
mild fatty infiltration of the liver | 0
managed conservatively | 0
treated with doxycycline 100 mg twice daily | 0
defervescence | 48
improved orientation | 48
weakness of both lower limbs (Grade 2/5) | 96
weakness progressed to upper limbs (Grade 2/5) | 96
absent deep tendon reflexes | 96
flexor plantar responses | 96
bladder incontinence | 96
no bowel incontinence | 96
breathing difficulty | 96
respiratory distress | 96
shifted to ICU | 96
single breath count 10 | 96
respiratory acidosis | 96
intubated | 96
mechanical ventilation | 96
MRI brain without any abnormality | 96
MRI cervical spine no abnormality | 96
motor sensory demyelinating polyneuropathy | 96
GBS | 96
CSF protein 146 | 96
CSF cell count 70 | 96
CSF lymphocytic predominance | 96
CSF sugar 71 mg/dL | 96
corresponding blood sugar 145 mg/dL | 96
intravenous immunoglobulin therapy 0.4 mg/kg/day | 96
tablet rifampicin 600 mg twice daily | 96
improvement in weakness of all four limbs | 144
improvement in respiratory parameters | 144
gradually weaned off ventilator | 144
extubated | 144
total duration of mechanical ventilation 10 days | 144
oral feeding started | 144
aggressive limb physiotherapy | 144
aggressive chest physiotherapy | 144
shifted out from ICU | 144
discharged from the hospital | 672
full neurological recovery | 672
total duration of hospital stay 4 weeks | 672
followed up regularly in outpatient department | 672
no functional disability | 672
