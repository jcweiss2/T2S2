38 years old| 0
female | 0
admitted to the hospital | 0
septic shock | 0
streptococcal necrotising fasciitis | 0
left chest wall | 0
amoxicilline | 0
clindamycine | 0
linezolid | 0
minor thoracic trauma | -48
playing sport | -48
infection spread to surface | -24
infection spread to pleura | -24
pneumothorax | -24
polymicrobial infection | 0
Stenotrophomonas maltophilia | 0
Citrobacter spp. | 0
Aspergillus spp. | 0
Mucor spp. | 0
refractory after 9 days of intensive treatment | 216
liposomal amphotericin B | 216
transferred to institution | 216
HBOT therapy | 216
Enterococcus faecium | 0
Enterobacter gallinarum | 0
Pseudomonas aeruginosa | 0
Citrobacter sedlakii | 0
Stenotrophomonas maltofilia | 0
Candida albicans | 0
Aspergillus fumigatus | 0
Aspergillus terreus | 0
mucormycosis | 264
Lichtheimia ramosa | 264
Rhizopus arrhizus | 264
cefepime | 264
ciprofloxacine | 264
sulfamethoxazole-trimethoprime | 264
metronidazole | 264
liposomal amphotericin B (67 days) | 264
pozaconazole (75 days) | 264
isavuconazole | 264
daily debridement surgery | 264
HBOT sessions | 264
vacuum therapy | 600
fungizone | 600
organ failures stabilised | 0
vasopressors weaning | 0
acute kidney injury | 0
continuous renal replacement therapy | 0
coagulopathy | 0
thrombocytopenia | 0
severe monocyte deactivation | 264
mHLA-DR < 5000 AB/C | 264
IFN-γ (100 mcg daily from day 11 to 21) | 264
increased mHLA-DR | 264
T lymphocyte PD-1 expression | 648
nivolumab (280 mg) | 648
IFN-γ on days 27, 28, and 31 | 648
PD-1 expression negative | 648
tissue culture negative for fungi | 672
blood PCR negative for fungi | 816
clinical status improved | 816
RRT weaning | 936
extubation | 1032
reconstructive surgery | 1248
skin grafting | 1248
left hospital | 3264
38 years old|0
female|0
admitted to the hospital|0
septic shock|0
streptococcal necrotising fasciitis|0
left chest wall|0
amoxicilline|0
clindamycine|0
linezolid|0
minor thoracic trauma|-48
playing sport|-48
infection spread to surface|-24
infection spread to pleura|-24
pneumothorax|-24
polymicrobial infection|0
Stenotrophomonas maltophilia|0
Citrobacter spp.|0
Aspergillus spp.|0
Mucor spp.|0
refractory after 9 days of intensive treatment|216
liposomal amphotericin B|216
transferred to institution|216
HBOT therapy|216
Enterococcus faecium|0
Enterobacter gallinarum|0
Pseudomonas aeruginosa|0
Citrobacter sedlakii|0
Stenotrophomonas maltofilia|0
Candida albicans|0
Aspergillus fumigatus|0
Aspergillus terreus|0
mucormycosis|264
Lichtheimia ramosa|264
Rhizopus arrhizus|264
cefepime|264
ciprofloxacine|264
sulfamethoxazole-trimethoprime|264
metronidazole|264
liposomal amphotericin B (67 days)|264
pozaconazole (75 days)|264
isavuconazole|264
daily debridement surgery|264
HBOT sessions|264
vacuum therapy|600
fungizone|600
organ failures stabilised|0
vasopressors weaning|0
acute kidney injury|0
continuous renal replacement therapy|0
coagulopathy|0
thrombocytopenia|0
severe monocyte deactivation|264
mHLA-DR < 5000 AB/C|264
IFN-γ (100 mcg daily from day 11 to 21)|264
increased mHLA-DR|264
T lymphocyte PD-1 expression|648
nivolumab (280 mg)|648
IFN-γ on days 27, 28, and 31|648
PD-1 expression negative|648
tissue culture negative for fungi|672
blood PCR negative for fungi|816
clinical status improved|816
RRT weaning|936
extubation|1032
reconstructive surgery|1248
skin grafting|1248
left hospital|3264
