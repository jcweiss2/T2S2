Here is the table of events and timestamps:

age | 65
sex | 0
admitted to the hospital | 0
history of shortness of breath | -4
fever | -4
cough | -4
fatigue | -4
oxygen saturation (SpO2) | -4
breath sounds reduced in the lower segments of the lungs | -4
nasopharyngeal SARS-CoV-2 RT-PCR test positive | -4
white cell count | -4
hemoglobin | -4
platelet count | -4
Westergren ESR | -4
interleukine 6 | -4
С-reactive protein | -4
ferritin | -4
D-dimer | -4
procalcitonin | -4
treated with dexamethason | -4
treated with heparin | -4
treated with tocilizumab | -4
treated with acetylcysteine | -4
treated with pantoprazole | -4
treated with nadroparin calcium | -4
oxygen supplementation | -4
chest CT scans | -4
bilateral peripheral ground-glass attenuation and patchy consolidation | -4
lung involvement 60%-70% | -4
positive for SARS-CoV-2 | -4
negative SARS-CoV-2 test result | -21
symptoms worsened | -21
increased temperature | -21
oxygen saturation (SpO2) decreased to 90% | -21
treated with linezolid | -21
treated with imipenem/cilastatin | -21
daily drainage volume | -21
pleural effusion with gas bubbles | -21
focal area of subpleural infiltration with a central cavity of destruction | -21
air layer up to 47 mm of anteroposterior thickness | -21
pleural effusion with 25 mm of anteroposterior depth | -21
air layer up to 19 mm of anteroposterior thickness | -21
multiple bilateral ground glass infiltrates | -21
pleural fluid analysis | -21
exudative lymphocytic-rich effusion | -21
no growth of acid-fast bacteria (AFB) | -21
Acinetobacter baumannii cultured | -21
Pseudomonas aeruginosa cultured | -21
Klebsiella pneumonia in urine culture | -21
needle thoracocentesis and new pleural drainage | -21
air and creamy purulent mass aspirated | -21
serofibrinous hemorrhagic fluid drawn daily | -21
chest CT showed air and pleural effusion in the right hemithorax | -21
diagnosis of pleural empyema | -21
transferred to the Surgical Department | -21
right pleural space irrigated with antiseptic solutions | -21
lung expansion by continuous vacuum aspiration technique | -21
encapsulated pleural effusion identified | -16
ultrasound-guided puncture of the effusion | -16
new drainage of the pleural cavity | -16
chest CT showed the presence of the encapsulated pleural effusion | -16
treated with colistimethatum natrium | -16
treated with imipenem/cilastatin | -16
discharged from the hospital | 24
oxygen saturation (SpO2) 97% on room air | 24
chest CT showed a small amount of fluid in the right pleural cavity | 24
lab test scores returned to normal range | 24
С-reactive protein 11.7 mg/l | 24
procalcitonin < 0.1 ng/ml | 24