12 years old | 0
female | 0
admitted to the emergency department | 0
complaining of anuria | 0
vomiting | 0
abdominal pain | 0
undergone severe Type III FGM | -2160
increasing pain during micturition | -2160
history of obstructed micturition | -2160
disrupted urinary stream | 0
splashing of very little urine | 0
malnourished | 0
tired | 0
in pain | 0
labia majora and minora amputated completely | -2160
fused labia minora remnant enclosing the vestibule | -2160
external urethral meatus and introitus covered entirely | -2160
anemic | 0
hemoglobin level of 5.9 g/dl | 0
creatinine 10.8 mg/dL | 0
urea 180 mg/dL | 0
leucocytes in urinalysis | 0
blood in urinalysis | 0
proteins in urinalysis | 0
urine culture showed growth of Escherichia Coli | 0
increased echogenicity in the bilateral renal parenchyma | 0
grade II renal parenchymal disease | 0
abdominal ascites | 0
hospitalized in the pediatric department | 0
obstructive nephropathy | 0
retention of urine | 0
bladder catheterization attempted | 0
impossible due to urethral meatus occluded and traumatized | 0
consultation with obstetrics and gynecology doctors | 0
decision for emergency defibrillation | 0
consent taken from the family | 0
emergency defibrillation surgery | 24
splitting the fused labia minora | 24
catheterization | 24
cut edges of the labia minora sutured together | 24
treatment at the pediatric intensive care units | 24
renal failure management started | 24
hemodialysis | 24
blood transfusion | 24
antibiotics | 24
condition deteriorating gradually | 48
lost her life due to sepsis | 72
sepsis resulted from chronic infection caused by FGM | 72