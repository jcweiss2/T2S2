66 years old | 0
female | 0
prior TIA | -120
urea cycle disorder | -8760
elevations of amino acids | -8760
genetic testing | -8760
OTC coding gene deletion | -8760
admitted to hospital | -240
confusion | -240
gait disturbance | -240
facial droop | -240
evaluation for stroke | -240
brain MRI | -240
brain toxicity | -240
encephalopathy | -240
increased ammonia level | -240
hallucinations | -48
worsening ataxia | -48
fall | -48
abdominal pain | -48
lower-extremity lymphedema | -48
elevated ammonia level | -48
hypoglycemia | -48
drop in hemoglobin | -48
hypotensive | 0
seizure | 0
Lorazepam | 0
normal saline bolus | 0
transferred to ICU | 0
blood pressure improvement | 0
albumin | 0
responsive | 0
Raviciti | 0
lactulose | 0
hyperammonemia | 0
vasopressors | 0
nosocomial pneumonia | 24
septic shock | 24
respiratory status worsening | 24
intubation | 24
vasopressor support | 24
ammonia levels fluctuation | 24
mental status fluctuation | 24
glucose levels fluctuation | 24
euglycemic state | 24
glucose fractioned solutions | 24
D5 | 24
D10 | 24
D20 | 24
normal saline | 24
persistent hypoglycemia | 24
HAHI syndrome | 24
genetic testing | 48
GLUD-1 gene mutation | 48
alpha-keto glutarate elevation | 48
ATP elevation | 48
insulin secretion | 48
hypoglycemia symptoms | 48
dizziness | 48
sweating | 48
confusion | 48
blurred vision | 48
balanced treatment | 72
dextrose 20 infusion | 72
Raviciti | 72
low-protein restricted diet | 72
mentation improvement | 72
registered dieticians | 72
metabolic disorders | 72
D20 infusion | 120
Raviciti | 120
low-protein restricted diet | 120
euglycemic level | 120
normal ammonia level | 120
discharged | 240