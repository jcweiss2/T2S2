67 years old | 0
female | 0
near-obstructing adenocarcinoma of the right colon | -120
laparoscopic-assisted extended right hemicolectomy | -120
discharged | -120
diffuse abdominal pain | -96
hematemesis | -96
subjective fevers | -96
free intraperitoneal fluid | -96
pneumoperitoneum | -96
broad spectrum antibiotics | -96
exploratory laparotomy | -96
anastomotic leak | -96
resection of anastomosis | -96
end ileostomy | -96
low grade tachycardia | -96
persistent obtundation | -24
extubation | -24
oxygen saturation above 95% | -24
apneic | -24
bag valve mask ventilation | -24
naloxone | -24
glycopyrrolate | -24
neostigmine | -24
profound respiratory acidosis | -24
pH of 7.03 | -24
PCO2 of 107 | -24
PaO2 of 375 | -24
re-intubation | -24
hypercapnic respiratory failure | -24
cerebral imaging | 0
acute cerebellar herniation | 0
diffuse cerebral edema | 0
decompressive external ventricular drain | 0
maximal medical therapy | 0
hypertonic saline | 0
head of bed elevation | 0
normotension | 0
normoglycemia | 0
levetiracetam | 0
seizure prophylaxis | 0
MRI | 0
PRES diagnosis | 0
vasogenic edema | 0
neurologic recovery | 240
discharged to rehabilitation facility | 240
ileostomy reversal | 720
complete resolution of neurological symptoms | 720
normalization of neuroimaging | 720