59 years old | 0
    male | 0
    non-obstructive hypertrophic cardiomyopathy | 0
    hospitalized | 0
    cardiac insufficiency | 0
    inotropic therapy | 0
    worsening of clinical picture | 0
    use of intra-aortic balloon | 0
    prioritized for cardiac transplantation | 0
    pre-transplant period | 0
    infectious complications | 0
    blood cultures | -48
    blood cultures | -24
    bicaval-bipulmonary heart transplantation | 0
    surgery | 24
    hemostasis | 24
    mechanical ventilation | 0
    vasoactive drugs | 0
    intra-aortic balloon | 0
    good clinical condition | 0
    mycophenolate mofetil | 0
    cyclosporine | 0
    prednisone |A 59-year-old male patient with non-obstructive hypertrophic cardiomyopathy was hospitalized to manage cardiac insufficiency with inotropic therapy. The worsening of his clinical picture required the use of an intra-aortic balloon, and he was prioritized for cardiac transplantation. During the pre-transplant period, the patient did not develop any infectious complications. Blood cultures collected 24 and 48 h before transplantation were negative.
    
    The patient underwent bicaval–bipulmonary heart transplantation, which required another surgery in the first 24 h to resolve hemostasis. He remained under mechanical ventilation with the use of vasoactive drugs and an intra-aortic balloon for 48 h, maintaining a good clinical condition. The immunosuppressive regimen included mycophenolate mofetil, cyclosporine and prednisone. On day 3 post-operation, a blood culture from the donor was positive for Gram-negative bacilli. As the donor was receiving piperacillin–tazobactam at the time of transplantation, the same drug was administered to the recipient. Although the recipient was clinically stable without signs of infection, blood cultures and surveillance cultures (from the groin and rectal areas) were collected. On day 5 post-operation, the final identification turned out ColR KPC-Kp.
    
    Blood cultures from the recipient were positive for ColR KPC-Kp on day 7 post-operation with the same sensitivity profile as the donor isolate. The surveillance cultures were negative. At this time, the recipient was afebrile and hemodynamically stable, presenting with 26,000 cells/mm3 leukocyte count and 6.5 mg/dL C-reactive protein (CRP) levels. Double-carbapenems (meropenem 2 g 8/8 h in a 4-h infusion combined with ertapenem 1 g/day, 1 h before one of the meropenem doses) and amikacin (15 mg/kg once a day) was started. The patient developed pericarditis on day 9 post-operation and required the drainage of 1000 mL of exudate; his pericardial fluid cultures were positive for ColR KPC-Kp. The patient underwent a surgical approach to clean the pericardium, requiring a repeated surgery eight days later; a sternum bone fragment collected at this time was positive for ColR KPC-Kp. On day 37 post-operation, he presented with worsening respiratory signs with chest computed tomography exhibiting consolidation with lung fluid levels suggestive of pulmonary cavitation due to necrosis (Fig. 1). This diagnosis was confirmed by histopathology of lung fragments obtained from lobectomy, in which a pulmonary abscess with liquefactive necrosis and necrotizing arteritis were noted. The patient developed septic shock, and antibiotic coverage was extended to linezolid and fluconazole while maintaining the initial treatment regimen for ColR KPC-Kp (double-carbapenem and amikacin). The patient progressed to multiple organ failure and died on day 50 post-transplantation.