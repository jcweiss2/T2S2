48 years old | 0
male | 0
admitted to the hospital | 0
pain | -2
distension of abdomen | -2
low-grade fever | -720
cough | -720
scanty expectoration | -720
weight loss | -720
anti-tubercular therapy | -720
bilateral upper zone opacities | -720
pulse rate 112/min | 0
blood pressure 134/86 mm of Hg | 0
respiratory rate 36/min | 0
temperature 100°F | 0
abdomen distended | 0
abdomen tender | 0
abdomen rigid | 0
abdomen guarding | 0
tenderness aggravated by movement | 0
tenderness aggravated by cough | 0
percussion note tympanitic | 0
vesicular breath sounds diminished intensity | 0
coarse crackles bilaterally | 0
hemoglobin 110 g/L | 0
total leukocyte count 11.2 × 10^9/L | 0
neutrophil 68% | 0
lymphocytes 27% | 0
polymorphonuclear leukocytosis | 0
liver enzymes mildly elevated | 0
aspartate transaminase 64 U/L | 0
alanine transaminase 78 U/L | 0
alkaline phosphatase 156 U/L | 0
random plasma glucose 98 mg/dL | 0
blood urea nitrogen 12 mmol/L | 0
creatinine 1.1 μmol/L | 0
sodium 134 mEq/L | 0
potassium 3.4 mEq/L | 0
serum amylase normal | 0
serum lipase normal | 0
urine examination normal | 0
HbSAg negative | 0
anti-hepatitis C virus negative | 0
HIV negative | 0
infiltrations in bilateral upper zones | -720
increased broncho vascular markings | -720
free gas under the diaphragm | 0
intraperitoneal gaseous distension | 0
intraperitoneal free fluids | 0
exploratory laparotomy | 2
purulent fluid | 2
perforations | 2
peritoneal lavage | 2
omentum fat | 2
pelvic drain | 2
mechanical ventilation | 2
piperacillin-tazobactam | 2
amikacin | 2
Gram-negative bacilli | 48
bipolar staining | 48
lactose fermenting pink colonies | 48
dry and wrinkled colonies | 96
ceftazidime | 120
amikacin | 120
B. pseudomallei | 144
imipenem | 144
doxycyclin | 144
T-piece ventilation | 216
oxygen | 216
T-piece removed | 288
oxygen saturation maintained | 288
imipenem stopped | 336
doxycyclin stopped | 336
cotrimoxazole | 336
discharged | 576
follow-up | 1296
no relapse | 1296