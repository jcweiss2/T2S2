62 years old | 0
    man | 0
    admitted to hospital | 0
    lumbar back pain | -168
    fever | -168
    chronic congestive heart failure | 0
    hypertension | 0
    diabetes mellitus | 0
    peripheral arterial disease | 0
    atrial fibrillation | 0
    hemodynamically stable | 0
    no acute signs of worsening cardiac function | 0
    no acute signs of worsening lung function | 0
    abdomen diffusely tender on palpation | 0
    no signs of peritoneal inflammation | 0
    non-contrast computed tomography scan | 0
    confluent mass of periaortic soft tissue | 0
    retroperitoneal fibrosis | 0
    aortic calcifications | 0
    urgent laboratory tests | 0
    12.280/mmc leukocytes | 0
    96% neutrophils | 0
    C-reactive protein of 225 mg/L | 0
    magnetic resonance imaging of dorsal and lumbar spine | 0
    no spondylodiscitis | 0
    transthoracic echocardiogram | 0
    no cardiac vegetations | 0
    intravenous meropenem | 0
    intravenous vancomycin | 0
    blood cultures positive for MSSA | 0
    treatment changed to intravenous cloxacillin | 0
    new onset syncope | 168
    shock | 168
    progressively worsening lumbar pain | 168
    repeat abdominal CT scan | 168
    retroperitoneal collection of blood | 168
    aortic rupture | 168
    left renal artery rupture | 168
    angiography confirmed CT findings | 168
    aortic balloon inflated above superior mesenteric artery | 168
    occluded vessel | 168
    endovascular aortic cuff placed at renal arteries | 168
    transferred to ICU | 168
    repeat abdominal and pelvis CT scan | 192
    small leak to right renal artery | 192
    patency of celiac trunk | 192
    patency of SMA | 192
    patency of right renal artery | 192
    patency of inferior mesenteric artery | 192
    operated on again | 288
    right colon ischemia | 288
    transverse colon ischemia | 288
    left colon ischemia | 288
    resection performed | 288
    repeat abdominal CT scan | 408
    no endoleak | 408
    patency of splachnic arteries except left renal | 408
    dependent on vasopressor | 0
    dependent on inotropic support | 0
    mechanical ventilation | 0
    hemodialysis | 0
    treated with vancomycin | 0
    treated with cloxacillin | 0
    persistence of MSSA bacteremia | 0
    patient expired | 408
    autopsy revealed mycotic thrombosed abdominal aneurysm | 408
    necrosis of left aortic wall | 408
    thrombosis of left renal artery | 408
    no aortic rupture | 408
    aortic wall infiltrated with neutrophils | 408
    gram positive cocci present | 408
    no endocardial vegetations | 408
    no valvular vegetations | 408
    no fibrotic tissue on peritoneum | 408
    multiple abscesses of peritoneal fat | 408
    bacterial invasion | 408
    yeast invasion | 408
    vascular invasion | 408