49 years old | 0
male | 0
admitted to the hospital | 0
chronic kidney disease | -23680
chronic glomerulonephritis | -23680
hypertension | -23680
hemodialysis | -23680
kidney transplant | -23680
antibody-mediated rejection | -23664
cytomegalovirus colitis | -23652
cyclosporin | -23680
ketoconazole | -23680
azathioprine | -23680
prednisone | -23680
lansoprazole | -23680
amlodipine | -23680
cough | -168
fever | -168
shortness of breath | -168
myalgia | -168
SARS-CoV-2 | -168
high-flow nasal oxygen | 0
fraction of inspired oxygen | 0
nasal prong oxygen | 0
immunosuppression | 0
anticoagulation | 0
enoxaparin | 0
corticosteroids | 0
increased prednisone | 0
chest X-ray | 0
bilateral diffuse infiltrates | 0
COVID-19 pneumonia | 0
creatinine | 0
urea | 0
potassium | 0
white cell count | 0
C-reactive protein | 0
D-dimer | 0
ferritin | 0
temperature spike | 48
urine cultures | 48
blood cultures | 48
carbapenem | 48
nosocomial sepsis | 48
noncontrast computed tomography | 72
abdomen | 72
chest | 72
pain over the graft kidney | 72
nephrology team | 72
ertapenem | 72
sodium polystyrene sulfonate | 72
hyperkalemia | 72
azathioprine discontinued | 72
hemodialysis | 120
refractory hyperkalemia | 120
metabolic acidosis | 120
sodium bicarbonate | 120
polyuric | 144
urine output | 144
cyclosporin level | 168
ketoconazole stopped | 168
cyclosporin increased | 168
graft kidney biopsy | 168
renal infarction | 168
graft loss | 168
discharge | 216
anticoagulation strategy | 216
kidney replacement therapy | 216
long-term anticoagulation | 216