72 years old | 0
    male | 0
    hypertension | 0
    atrial fibrillation | 0
    alcoholic liver cirrhosis | 0
    metastatic urothelial carcinoma | 0
    presented to the hospital for evaluation of rash | 0
    rash developed shortly after day 8 infusion | -168
    scheduled to receive enfortumab vedotin on days 1, 8, and 15 | -168
    tolerated day 1 well | -168
    day 8 infusion | -168
    erythematous rash with skin sloughing on <20% of body | -168
    admitted to M.D. Anderson Cancer Center | -144
    rash progressed | -144
    transferred to burn intensive care unit on day 12 | -144
    hemodynamically stable on admission | 0
    tense bullae on background of erythema on bilateral axillae | 0
    tense bullae on background of erythema on back | 0
    tense bullae on background of erythema on genitalia | 0
    tense bullae on background of erythema on posterior aspect of bilateral thighs | 0
    tense bullae on background of erythema on bilateral heels | 0
    single blister on posterior aspect of oral cavity | 0
    concern for Stevens-Johnson syndrome/TEN | 0
    SCORTEN score 7 | 0
    ABCD-10 score 5 | 0
    medication review | 0
    acetaminophen | 0
    acyclovir | 0
    metoprolol | 0
    gabapentin | 0
    no recent dose changes | 0
    no recent antiepileptics | 0
    no recent antibiotics | 0
    recent initiation of enfortumab vedotin | -168
    rapid-onset development of rash | -168
    enfortumab vedotin discontinued | 0
    started on topical steroid | 0
    biopsy performed | 0
    interface dermatitis with full-thickness epidermal necrosis | 0
    consistent with SJS/TEN overlap | 0
    oliguria developed overnight | 24
    urine microscopy revealed muddy brown casts | 24
    acute kidney injury secondary to acute tubular necrosis | 24
    started on continuous renal replacement therapy | 24
    rash progressed to involve >30% of skin | 24
    diagnosed with TEN | 24
    systemic steroids contraindicated | 24
    condition deteriorated | 24
    discussed treatment options | 24
    considered intravenous immunoglobulin | 24
    considered cyclosporine | 24
    considered etanercept | 24
    continued on supportive therapy | 24
    empiric vancomycin/meropenem | 24
    day 3 of hospitalization | 72
    SCORTEN remained at 7 | 72
    hypotension did not resolve | 72
    started on norepinephrine | 72
    started on vasopressin | 72
    laboratory evidence of hyperbilirubinemia | 72
    increased international normalized ratio | 72
    MELD score increased to 40 | 72
    multiorgan failure | 72
    septic shock | 72
    end-of-life measures discussed | 72
    died 20 days after admission | 480
    <|eot_id|>
