29 years old | 0
male | 0
admitted to the hospital | 0
asthma | 0
previous gunshot wound | 0
obesity | 0
tobacco use | 0
worked at auto-parts manufacturing unit | 0
dyspnea | -72
cough | -72
fatigue | -72
myalgias | -72
febrile | 0
tachycardic | 0
tachypneic | 0
supplemental oxygen | 0
ill appearance | 0
high work of breathing | 0
productive cough | 0
lymphopenia | 0
thrombocytopenia | 0
unremarkable chest radiograph | 0
transferred to ICU | 0
high suspicion for COVID-19 | 0
SARS-CoV-2 testing | 0
nasopharyngeal swab | 0
chest CT not performed | 0
required higher flow rates on non-rebreather mask | 72
persistent fevers | 96
tachypnea | 96
new consolidative changes in right middle and lower lung zones | 96
broad-spectrum antibiotics | 96
hydroxychloroquine | 96
mechanical ventilation | 96
extensive consolidative infiltrates bilaterally | 192
PaO2/FiO2 ratio of 59 | 192
severe ARDS | 192
SARS-CoV-2 positive | 192
septic shock | 192
vasopressor support | 192
IL-6 of 46 pg/mL | 192
cytokine release syndrome | 192
tocilizumab 400 mg | 192
extensive acute DVTs in left upper extremity | 240
d-dimer levels over 10 µg/mL | 240
enoxaparin increased to therapeutic dose | 240
fevers not abated | 240
cooling | 240
neuromuscular blockade | 240
deep sedation | 240
ARDS strategies | 240
low tidal volumes | 240
proning | 240
recruitment maneuvers | 240
diuretics | 240
nitric oxide | 240
vitamin C | 240
high plateau pressures | 240
consideration of ECMO transfer | 240
left-sided tension pneumothorax | 408
chest tube draining 700 mL serosanguineous fluid | 408
persistent air leaks | 408
desaturation | 408
family discussion | 408
DNR | 408
asystole | 480
death | 480
obesity |@0
tobacco use |@0
worked at auto-parts manufacturing unit |@0
dyspnea |@-72
cough |@-72
fatigue |@-72
myalgias |@-72
febrile |@0
tachycardic |@0
tachypneic |@0
supplemental oxygen |@0
ill appearance |@0
high work of breathing |@0
productive cough |@0
lymphopenia |@0
thrombocytopenia |@0
unremarkable chest radiograph |@0
transferred to ICU |@0
high suspicion for COVID-19 |@0
SARS-CoV-2 testing |@0
nasopharyngeal swab |@0
chest CT not performed |@0
required higher flow rates on non-rebreather mask |@72
persistent fevers |@96
tachypnea |@96
new consolidative changes in right middle and lower lung zones |@96
broad-spectrum antibiotics |@96
hydroxychloroquine |@96
mechanical ventilation |@96
extensive consolidative infiltrates bilaterally |@192
PaO2/FiO2 ratio of 59 |@192
severe ARDS |@192
SARS-CoV-2 positive |@192
septic shock |@192
vasopressor support |@192
IL-6 of 46 pg/mL |@192
cytokine release syndrome |@192
tocilizumab 400 mg |@192
extensive acute DVTs in left upper extremity |@240
d-dimer levels over 10 µg/mL |@240
enoxaparin increased to therapeutic dose |@240
fevers not abated |@240
cooling |@240
neuromuscular blockade |@240
deep sedation |@240
ARDS strategies |@240
low tidal volumes |@240
proning |@240
recruitment maneuvers |@240
diuretics |@240
nitric oxide |@240
vitamin C |@240
high plateau pressures |@240
consideration of ECMO transfer |@240
left-sided tension pneumothorax |@408
chest tube draining 700 mL serosanguineous fluid |@408
persistent air leaks |@408
desaturation |@408
family discussion |@408
DNR |@408
asystole |@480
death |@480
