50 years old | 0
female | 0
presented | 0
fever | -168
abdominal pain | -168
loose stools | -168
dry cough | -336
symptomatic treatment | -336
no vomiting | 0
no dyspnoea | 0
no sputum production | 0
no haemoptysis | 0
no previous history of obstructive airway disease | 0
no antitubercular treatment |==0
type 2 diabetes mellitus | -17520
hypertension | -17520
hypothyroidism | -17520
regular medicines | -17520
thyroid surgery | -157680
multinodular goitre | -157680
surgical site infection | -157848
tracheal involvement | -157848
on and off dry cough | -70080
cough suppressants | -70080
antibiotics | -70080
symptoms recurrence | -70080
moderately built | 0
weight 62 kg | 0
afebrile | 0
blood pressure 80/50 mmHg | 0
pulse rate 110/min |
