12 years old | 0
female | 0
admitted to the hospital | 0
fever | -336
joint swelling | -336
joint pain | -336
hair lice | -336
scratch marks on scalp | -336
bilateral pleural effusion | 0
ejection systolic murmur | 0
tender hepatomegaly | 0
multiple joint swelling | 0
multiple joint redness | 0
multiple joint tenderness | 0
increased WBC count | 0
lymphocytes 0.9×10^9 cells/l | 0
granulocytes 4.5×10^9 cells/l | 0
monocytes 0.2×10^9 cells/l | 0
reticulocytes 28×10^9 cells/l | 0
thrombocytopenia | 0
anemia | 0
hyponatremia | 0
hyperkalemia | 0
hypoglycemia | 0
elevated serum urea | 0
elevated serum creatinine | 0
elevated LDH | 0
elevated AST | 0
elevated ALT | 0
elevated ALP | 0
hypoalbuminemia | 0
elevated GGT | 0
elevated CK | 0
hyperbilirubinemia | 0
serum osmolality 289 mOsm/kg | 0
urine osmolality 647 mOsm/kg | 0
INR 1.2 | 0
prothrombin time 14 | 0
activated partial thromboplastin time 36 | 0
anti-hepatitis B surface antigen positive | 0
chest X-ray showed bilateral pleural effusion | 0
chest X-ray showed widened mediastinum | 0
ECG showed sinus tachycardia | 0
ECG showed diffuse ST-segment elevation | 0
ECG showed generalized T-wave inversion | 0
transthoracic echocardiogram showed moderate pericardial effusion | 0
blood cultures obtained | 0
sputum cultures obtained | 0
urine cultures obtained | 0
ceftazidime started | 0
flucloxacillin started | 0
right chest tube thoracostomy inserted | 0
pleural fluid analysis | 0
Gram-positive cocci in clusters seen on Gram stain | 0
hair shaved | 0
anti-lice shampoo started | 0
sputum microscopy negative for acid-fast bacilli | 0
mycobacterium tuberculosis culture sent | 0
polymerase chain reaction test sent | 0
intubated | 24
mechanical ventilation started | 24
antibiotics changed to meropenem | 24
dopamine infusion started | 24
norepinephrine infusion started | 24
air leak from right chest tube observed | 24
echocardiography-guided pericardiocentesis performed | 24
pericardial fluid analysis | 24
pericardial fluid showed proteins 42 g/l | 24
pericardial fluid showed albumin 27 g/l | 24
pericardial fluid showed Gram-positive cocci in clusters | 24
chest X-ray showed right minimal hydropneumothorax | 24
ultrasound examination of abdomen showed perinephric collections | 24
ultrasound examination of abdomen showed subhepatic collections | 24
ultrasound examination of abdomen showed free fluid in abdomen and pelvis | 24
methicillin-sensitive Staphylococcus aureus cultured from sputum | 24
methicillin-sensitive Staphylococcus aureus cultured from blood | 24
methicillin-sensitive Staphylococcus aureus cultured from pleural fluid | 24
methicillin-sensitive Staphylococcus aureus cultured from pericardial aspirate | 24
urine cultures negative | 24
rheumatoid factor levels slightly elevated | 24
cytomegalovirus IgM antibodies negative | 24
cytomegalovirus IgG titer 1/21,000 IU/L | 24
air leak through pericardial pig-tail catheter observed | 72
broncho-pericardial or broncho-pleuropericardial fistula suspected | 72
pig-tail catheter clamped | 72
BP decreased to 80/50 mmHg | 72
HR increased to 120 beats/min | 72
pig-tail catheter de-clamped | 72
BP returned to baseline | 72
HR returned to baseline | 72
CT of chest showed pneumopericardium | 72
CT of chest showed hydropneumothorax | 72
CT fistulogram confirmed communication between right pleural space and pericardium | 72
conservative management recommended | 72
abdominal collections aspirated laparoscopically | 96
disseminated intravascular coagulation developed | 216
bleeding from everywhere | 216
died of multi-organ failure | 264
autopsy refused | 264