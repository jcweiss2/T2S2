13 years old | 0
male | 0
scheduled for elective insertion of a continuous ambulatory peritoneal dialysis (CAPD) catheter | 0
admission height 135 cm | 0
admission weight 31 kg | 0
born at 40 weeks | -105120
normal vaginal delivery | -105120
admitted to the neonatal intensive care unit | -105120
sepsis | -105120
mitochondrial disease diagnosed | -132192
Joubert syndrome diagnosed | -132192
hemodialysis started | -26208
end-stage renal disease | -26208
hospitalized with intracranial hemorrhage | -17520
high blood pressure | -17520
admitted for uncontrolled hypertension | -8760
change in the permanent catheter | -8760
hyperkalemia-induced cardiac arrest | -8760
cardiopulmonary resuscitation (CPR) | -8760
spontaneous circulation returned | -8760
transferred to the intensive care unit (ICU) | -8760
post-CPR care received for 2 weeks | -8760
hospitalized and discharged repeatedly due to heart, lung, and kidney problems | 0
regular hemodialysis | 0
hemoglobin level continued to fall | 0
blood pressure continued to fall | 0
scheduled to switch to peritoneal dialysis | 0
stuporous mental status | 0
Glasgow coma scale (GCS) score 11 | 0
-ridden | 0
percutaneous endoscopic gastrostomy tube inserted | 0
hypotension managed by norepinephrine infusion | 0
mean blood pressure (MBP) 90–106 mmHg | 0
heart rate (HR) 95–107 beats/min | 0
shallow breathing | 0
100% oxygen saturation maintained on room air | 0
no previous surgery | 0
small jaw | 0
slightly protruding mouth | 0
short neck | 0
reduced cervical mobility | 0
poor mouth opening | 0
rigidity of jaw | 0
blood sugar 132 mg/dl | 0
operating room NIBP 120/90 mmHg | 0
operating room HR 105 beats/min | 0
norepinephrine infusion 0.07 µg/kg/min | 0
invasive blood pressure monitoring not performed | 0
left radial artery cannulation prepared | 0
train-of-four (TOF) stimulation monitored | 0
bispectral index (BIS) 71 | 0
anesthesia started with propofol | 0
remifentanil | 0
rocuronium | 0
preoxygenation | 0
propofol infusion 77–102 µg/kg/min | 0
remifentanil infusion 0.05–0.1 µg/kg/min | 0
BIS maintained at 40–60 | 0
palate not malformed | 0
tongue not protruding | 0
mask ventilation well maintained | 0
I-gel insertion attempted | 0
air leak | 0
insufficient tidal volume | 0
I-gel removed | 0
trachea secured with endotracheal tube (ETT) | 0
Cormack-Lehane grade 1 | 0
pilot balloon inflated | 0
cuff pressure 18 cmH2O | 0
decreased lung sounds on left side | 0
coarse breath sounds over both lower lung fields | 0
ETT fixed at 15 cm | 0
mechanical ventilation settings | 0
50:50 air/oxygen mixture | 0
tidal volume 6–8 ml/kg | 0
respiratory rate 16–18 breaths/min | 0
maximum peak airway pressure 11–14 cmH2O | 0
inspiratory/expiratory time ratio 1:2 | 0
end-tidal carbon dioxide 35–39 mmHg | 0
oxygen saturation 100% | 0
operation duration 45 min | 0
MBP 73–103 mmHg | 0
HR 105–130 beats/min | 0
norepinephrine infusion 0.03–0.07 µg/kg/min | 0
TOF count 1–2 | 0
no additional muscle relaxants | 0
no additional opioids | 0
spontaneous breathing returned | 0
BIS 73 | 0
TOF ratio 76% | 0
respiration rate < 10 times/min | 0
midazolam injected | 0
transferred to SICU with ETT | 0
stuporous mental state (GCS score 6) | 24
ventilator applied | 24
synchronized intermittent mandatory ventilation mode | 24
FiO2 0.25 | 24
tidal volume 6 ml/kg | 24
respiratory rate 20 breaths/min | 24
pressure support 13 cmH2O | 24
MBP 105–111 mmHg | 24
HR 124–137 beats/min | 24
norepinephrine infusion 0.07 µg/kg/min | 24
trachea extubated | 24
no irregular respiratory patterns observed | 24
100% oxygen saturation with 2-L nasal cannula | 24
venous pH 7.30 | 24
PCO2 53 mmHg | 24
PO2 47 mmHg | 24
base excess 0.3 mmol/L | 24
SO2 78% | 24
glucose 130 mg/L | 24
lactate 0.3 mmol/L | 24
13 years old|0
male|0
scheduled for elective insertion of a continuous ambulatory peritoneal dialysis (CAPD) catheter|0
admission height 135 cm|0
admission weight 31 kg|0
born at 40 weeks|-105120
normal vaginal delivery|-105120
admitted to the neonatal intensive care unit|-105120
sepsis|-105120
mitochondrial disease diagnosed|-132192
Joubert syndrome diagnosed|-132192
hemodialysis started|-26208
end-stage renal disease|-26208
hospitalized with intracranial hemorrhage|-17520
high blood pressure|-17520
admitted for uncontrolled hypertension|-8760
change in the permanent catheter|-8760
hyperkalemia-induced cardiac arrest|-8760
cardiopulmonary resuscitation (CPR)|-8760
spontaneous circulation returned|-8760
transferred to the intensive care unit (ICU)|" -8760
post-CPR care received for 2 weeks|-8760
hospitalized and discharged repeatedly due to heart, lung, and kidney problems|0
regular hemodialysis|0
hemoglobin level continued to fall|0
blood pressure continued to fall|0
scheduled to switch to peritoneal dialysis|0
stuporous mental status|0
Glasgow coma scale (GCS) score 11|0
bed-ridden|0
percutaneous endoscopic gastrostomy tube inserted|0
hypotension managed by norepinephrine infusion|0
mean blood pressure (MBP) 90–106 mmHg|0
heart rate (HR) 95–107 beats/min|0
shallow breathing|0
100% oxygen saturation maintained on room air|0
no previous surgery|0
small jaw|0
slightly protruding mouth|0
short neck|0
reduced cervical mobility|0
poor mouth opening|0
rigidity of jaw|0
blood sugar 132 mg/dl|0
operating room NIBP 120/90 mmHg|0
operating room HR 105 beats/min|0
norepinephrine infusion 0.07 µg/kg/min|0
invasive blood pressure monitoring not performed|0
left radial artery cannulation prepared|0
train-of-four (TOF) stimulation monitored|0
bispectral index (BIS) 71|0
anesthesia started with propofol|0
remifentanil|0
rocuronium|0
preoxygenation|0
propofol infusion 77–102 µg/kg/min|0
remifentanil infusion 0.05–0.1 µg/kg/min|0
BIS maintained at 40–60|0
palate not malformed|0
tongue not protruding|0
mask ventilation well maintained|0
I-gel insertion attempted|0
air leak|0
insufficient tidal volume|0
I-gel removed|0
trachea secured with endotracheal tube (ETT)|0
Cormack-Lehane grade 1|0
pilot balloon inflated|0
cuff pressure 18 cmH2O|0
decreased lung sounds on left side|0
coarse breath sounds over both lower lung fields|0
ETT fixed at 15 cm|0
mechanical ventilation settings|0
50:50 air/oxygen mixture|0
tidal volume 6–8 ml/kg|0
respiratory rate 16–18 breaths/min|0
maximum peak airway pressure 11–14 cmH2O|0
inspiratory/expiratory time ratio 1:2|0
end-tidal carbon dioxide 35–39 mmHg|0
oxygen saturation 100%|0
operation duration 45 min|0
MBP 73–103 mmHg|0
HR 105–130 beats/min|0
norepinephrine infusion 0.03–0.07 µg/kg/min|0
TOF count 1–2|0
no additional muscle relaxants|0
no additional opioids|0
spontaneous breathing returned|0
BIS 73|0
TOF ratio 76%|0
respiration rate < 10 times/min|0
midazolam injected|0
transferred to SICU with ETT|0
stuporous mental state (GCS score 6)|24
ventilator applied|24
synchronized intermittent mandatory ventilation mode|24
FiO2 0.25|24
tidal volume 6 ml/kg|24
respiratory rate 20 breaths/min|24
pressure support 13 cmH2O|24
MBP 105–111 mmHg|24
HR 124–137 beats/min|24
norepinephrine infusion 0.07 µg/kg/min|24
trachea extubated|24
no irregular respiratory patterns observed|24
100% oxygen saturation with 2-L nasal cannula|24
venous pH 7.30|24
PCO2 53 mmHg|24
PO2 47 mmHg|24
base excess 0.3 mmol/L|24
SO2 78%|24
glucose 130 mg/L|24
lactate 0.3 mmol/L|24
