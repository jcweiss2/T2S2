69 years old | 0
    male | 0
    diabetes mellitus | 0
    hypertension | 0
    56 pack-year smoking | 0
    abdominal distension | 0
    abdominal pain | 0
    severe diffuse abdominal tenderness | 0
    rebound | 0
    guarding | 0
    peritonitis | 0
    white blood cell count 9.4 × 10^9 cells/L | 0
    hemoglobin 10.9 g/dL | 0
    platelets 370 × 10^9 cells/L | 0
    creatinine 1.29 mg/dL | 0
    thickening of the sigmoid colon | 0
    pneumoperitoneum | 0
    intraperitoneal free fluid | 0
    multifocal liver lesions | 0
    peritoneal implants | 0
    omental implants | 0
    metastatic perforated sigmoid carcinoma | 0
    exploratory laparotomy | 0
    perforated sigmoid | 0
    multiple liver lesions | 0
    omental lesions | 0
    sigmoidectomy | 0
    end colostomy | 0
    partial omentectomy | 0
    wedge resection of liver segment III | 0
    postoperative care | 0
    poorly differentiated squamous cell carcinoma | 0
    immunohistochemical staining primary pulmonary source | 0
    tumor cells positive CK5/6 | 0
    tumor cells positive p40 | 0
    tumor cells negative CK7 | 0
    tumor cells negative CK20 | 0
    tumor cells negative villin | 0
    tumor cells negative TTF1 | 0
    right perihilar mass | 0
    obstruction of right upper and middle lobe bronchi | 0
    encasement of right pulmonary artery branches | 0
    extensive bulky mediastinal lymphadenopathy | 0
    primary lung cancer | 0
    peritonitis secondary to perforated sigmoid mass | 0
    metastatic right lung squamous cell non-small cell lung cancer | 0
    acute abdominal symptoms as first manifestation of metastatic lung cancer | 0
    obstructive bronchopneumonia | 0