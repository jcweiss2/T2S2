17 years old | 0
male | 0
admitted to the intensive care unit | 0
fever | -48
diarrhea | -48
vomiting | -48
syncope | -48
pale | 0
febrile | 0
icteric | 0
tachycardic |)
hypotensive | 0
methicillin-sensitive Staphylococcus aureus blood cultures | 0
intravenous fluids | 0
dopamine 5 μg/kg/min | 0
intravenous vancomycin 1g every 12h | 0
rifampicin 300mg every 8h | 0
gentamicin 62mg every 12h | 0
vancomycin stopped | 0
intravenous oxacillin 2g every 4h | 0
right ventricular pressure normal | 0
right ventricular pressure increased to near-systemic | 48
stent precluding visualization of Melody valve leaflets | 0
cardiac magnetic resonance imaging no perivalvular abscess | 0
computed tomography chest multiple cavitary nodules | 0
septic emboli | 0
condition stabilized | 48
discharged from intensive care unit | 48
gentamicin stopped | 336
oxacillin treatment | 1008
rifampicin treatment | 1008
elective scheduled for Melody valve explantation | 1008
inflammation around calcified homograft | 1008
Melody valve infected | 1008
thickened valve leaflets | 1008
adhered valve leaflet | 1008
homograft explanted | 1008
Melody valve explanted | 1008
pulmonary homograft replacement | 1008
acute inflammatory infiltrate | 1008
granulation tissue | 1008
acute endocarditis | 1008
postoperative course uneventful | 1008
6 months follow-up well | 4032
complete transposition of the great arteries | -87600
ventricular septal defect | -87600
pulmonary stenosis | -87600
Rastelli repair | -87600
16mm pulmonary homograft | -87600
conduit replacement | -72240
20mm aortic homograft | -72240
balloon dilated | -52560
transcatheter Melody valve placed | -52560
minimal gradient across conduit | -43800
no more than mild regurgitation | -43800
history of prior endocarditis | -52560
male gender | -87600
previous endocarditis | -52560
prior stent implantations in RVOT | -52560
altered RVOT anatomy | -52560
stopped antiplatelet therapy | -52560
