27 years old | 0
    woman | 0
    gravida 2 para 0 | 0
    unremarkable medical history | 0
    unremarkable family history | 0
    admitted at 30 weeks and 3 days of pregnancy | 0
    abdominal pain | 0
    fever | 0
    body temperature 38.9°C | 0
    blood pressure 110/70 mmHg | 0
    heart rate 115 beats per minute | 0
    marked splenomegaly | 0
    no swelling of superficial lymph nodes | 0
    no tumor mass indicative of lymphoma | 0
    hemoglobin 7.9 g/dL | 0
    absolute neutrophil count 0.92 × 10^9/L | 0
    platelet count 25 × 10^9/L | 0
    elevated alanine aminotransferase 72 U/L | 0
    elevated aspartate aminotransferase 463 U/L | 0
    elevated lactate dehydrogenase 1799 U/L | 0
    elevated C-reactive protein 19.5 mg/dL | 0
    hypofibrinogenemia 0.94 g/L | 0
    elevated serum ferritin 438,600 ng/mL | 0
    prolonged prothrombin time (INR 1.90) | 0
    elevated fibrinogen degradation product 48.7 μg/mL | 0
    splenic swelling 9.8 cm thick | 0
    negative viral serology for HIV | 0
    negative viral serology for cytomegalovirus | 0
    negative viral serology for hepatitis B | 0
    negative viral serology for hepatitis C | 0
    no relief of presenting symptoms | 0
    alanine aminotransferase elevated to 163 U/L | 24
    aspartate aminotransferase elevated to 825 U/L | 24
    deteriorating general status | 24
    fetal distress | 24
    emergency cesarean section | 24
    1750 g male infant delivered | 24
    Apgar scores 5 to 8 points | 24
    neonatal respiratory distress syndrome | 24
    no macroscopic placental abnormalities | 24
    postoperation decline | 24
    disseminated intravascular coagulation | 24
    transfusion of 2 units packed red blood cells | 24
    transfusion of 2 units fresh frozen plasma | 0
    hemoglobin dropped to 5.7 g/dL | 24
    pink-tainted drainage fluid | 24
    spleen thickness 6.3 cm | 24
    probable postoperative abdominal hemorrhage | 24
    explorative laparotomy | 24
    ruptured spleen found | 24
    splenectomy performed | 24
    no improvement in condition | 24
    degrading liver function | 24
    acute respiratory distress | 24
    sustained kidney injury | 24
    transferred to intensive care unit | 24
    PiCCO monitor | 24
    CRRT | 24
    ventilator-assisted breathing | 24
    multiple blood products transfused | 24
    persistent cytopenia | 24
    persistent coagulopathy | 24
    deteriorating condition | 24
    bone marrow biopsy showing hemophagocytosis | 24
    atypical lymphoid cells | 24
    no abnormal clone cells in peripheral blood | 24
    no PNH clones in red and white blood cells | 24
    abnormal NK cells 3.57% | 24
    CD7 and cytoplasin attenuated expression | 24
    no expression of CD16 | 24
    no expression of CD11b | 24
    no expression of CD8 | 24
    no expression of CD57 | 24
    Ki67 positive ratio 28.8% | 24
    EBV serology positive | 24
    EBV DNA titer >1.0 × 10^7 | 24
    splenic rupture evidence | 24
    splenic corpuscle atrophy | 24
    splenic pulp hemophagocytosis | 24
    diffuse lymphoid cell infiltration | 24
    T cells infiltration | 24
    immunohistochemical staining CD56(+) | 24
    GrB(+) | 24
    TIA-1(+) | 24
    CD2(+) | 24
    CD3(part+) | 24
    CD5(−) | 24
    CD7(+) | 24
    CD43(+) | 24
    CD4(−) | 24
    CD8(−) | 24
    TdT(−) | 24
    CD20(−) | 24
    CD79α(−) | 24
    PAX-5(−) | 24
    CD34(−) | 24
    CD117(−) | 24
    MPO(−) | 24
    CD99(−) | 24
    CD123(−) | 24
    LCA(+) | 24
    CD68(−) | 24
    CD163(−) | 24
    Mum-1(−) | 24
    κ(−) | 24
    λ(−) | 24
    Ki-67(40%) | 24
    EBER CISH (+) | 24
    diagnosed invasive NK/T-cell lymphoma | 24
    diagnosed HLH | 24
    immunosuppressive therapy with dexamethasone | 24
    etoposide | 24
    rituximab | 24
    clinical symptoms deteriorated | 24
    died on 18th day postoperation | 432
    multiorgan failure | 432