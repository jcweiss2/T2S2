54 years old | 0
female | 0
HIV infection | -7200
admitted to the hospital | 0
complaints of pain over the right hip | 0
inability to bear weight on the right lower limb | 0
trivial fall | -1
tenderness over the right hip | 0
shortening of the right lower limb | 0
restricted range of motion | 0
fractured neck of the right femur | 0
azotemia | 0
hypokalemia | 0
anemia | 0
glycosuria | 0
proteinuria | 0
raised serum alkaline phosphatase level | 0
normal anion gap metabolic acidosis | 0
oral potassium supplementation | 0
modification of ART | 0
abacavir | 0
lamivudine | 0
efavirenz | 0
hemiarthroplasty | 0
urine routine and microscopic examination | 0
glucose 3+ | 0
protein 1+ | 0
few red blood cells | 0
no evidence of any crystals | 0
diagnosis of renal Fanconi syndrome | 0
hypokalemia | 0
hypophosphatemia | 0
glycosuria | 0
proteinuria | 0
hyperchloremic metabolic acidosis | 0
raised alkaline phosphatase levels | 0
serum 1,25-dihydroxyvitamin D level | 0
ultrasonography of the abdomen | 24
gross dilatation of the right kidney's pelvicalyceal system | 24
multiple calculi involving both the kidneys | 24
non-contrast computed tomographic imaging | 24
findings of USG were confirmed | 24
right kidney measured 9.8 cm | 24
normal contour and attenuation pattern | 24
four calculi noted in the right kidney's lower polar region | 24
largest measuring 2.1 cm × 1.6 cm | 24
few air pockets noted in the lower pole calyces | 24
emphysematous pyelitis | 24
6-mm calculus noted in the proximal right ureter | 24
causing upstream hydroureteronephrosis | 24
left kidney measured 8.3 cm | 24
normal contour and attenuation pattern | 24
calculus measuring 3 mm noted in the lower polar calyx of the right kidney | 24
cystopanendoscopy | 48
right double “J” stenting | 48
tachycardia | 72
tachypnea | 72
hypotension | 72
clinical diagnosis of pulmonary thromboembolism | 72
unfractionated heparin | 72
neutrophilic leucocytosis | 78
worsening azotemia | 78
arterial blood gas analysis showed severe metabolic acidosis | 78
urine culture had grown Escherichia coli | 78
Enterobacter aerogenes | 78
sensitive to ciprofloxacin | 78
piperacillin plus tazobactam | 78
culture-sensitive injectable antibiotics | 78
renal-modified doses | 78
bicarbonate infusion | 78
patient's condition improved | 150
extubated | 150
serum creatinine gradually improved | 150
discharged | 240
follow up after 1 month | 720