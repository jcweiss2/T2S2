46 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
ulcerative colitis | 0 | 0 | Factual
malaise | -72 | 0 | Factual
fever | -72 | 0 | Factual
loss of appetite | -72 | 0 | Factual
admitted to the hospital | 0 | 0 | Factual
blood pressure 124/46 mmHg | 0 | 0 | Factual
heart rate 122 beats per min | 0 | 0 | Factual
SpO2 98% | 0 | 0 | Factual
respiratory rate 16/min | 0 | 0 | Factual
body temperature 40.2°C | 0 | 0 | Factual
chills | 0 | 0 | Factual
nausea | 0 | 0 | Factual
cardiac arrest | 0 | 0 | Factual
chest compression | 0 | 0 | Factual
tracheal intubation | 0 | 0 | Factual
ventricular fibrillation | 0 | 0 | Factual
defibrillation | 0 | 0 | Factual
adrenaline administration | 0 | 0 | Factual
Brugada syndrome | 0 | 0 | Factual
coved-type ST elevation | 0 | 0 | Factual
hypercalcemia | 0 | 0 | Factual
serum calcium 14.8 mg/dL | 0 | 0 | Factual
hypotension | 0 | 24 | Factual
septic shock | 0 | 24 | Possible
ulcerative colitis exacerbation | 0 | 24 | Possible
tazobactam-piperacillin administration | 0 | 168 | Factual
vasopressors administration | 0 | 168 | Factual
extubation | 48 | 48 | Factual
fever reoccurred | 120 | 120 | Factual
liver abscess | 120 | 120 | Factual
meropenem administration | 120 | 504 | Factual
vancomycin administration | 120 | 504 | Factual
puncture drainage | 120 | 504 | Factual
infection controlled | 504 | 504 | Factual
pilsicainide test | 720 | 720 | Factual
implantable cardioverter defibrillator implantation | 720 | 720 | Factual
discharged | 720 | 720 | Factual
family history of sudden death | 0 | 0 | Factual
high parathyroid hormone levels | 720 | 720 | Factual
abnormal uptake in the anterior mediastinum | 720 | 720 | Factual
tumor resection | 720 | 720 | Factual
ectopic parathyroid adenoma | 720 | 720 | Factual
nonfunctional pituitary adenoma | 720 | 720 | Factual
nonfunctional adrenal tumor | 720 | 720 | Factual
multiple endocrine neoplasia type 1 | 720 | 720 | Factual