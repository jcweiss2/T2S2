69 years old | 0
female | 0
admitted to the senior behavioral health unit | 0
history of resected bifrontal meningioma | -672
breast cancer | -672
hypothyroidism | -672
pembrolizumab infusion | -48
altered mental status | -48
acute aphasia | -48
recurrent right facial twitching | -48
magnetic resonance imaging (MRI) brain | -48
chronic bifrontal encephalomalacia | -48
no acute ischemia on MRI brain | -48
continuous video EEG | -48
left frontal status epilepticus | -48
seizures treated with intravenous mid-azolam | -48
seizures treated with levetiracetam | -48
seizures treated with fosphenytoin | -48
seizures treated with valproic acid | -48
septic shock | -336
right lower lobe pneumonia | -336
vasopressor support | -336
mechanical ventilation | -336
lethargic | -336
cerebral spinal fluid (CSF) evaluation | -168
antiepileptic regimen tapered | -168
levetiracetam 500 mg twice daily | -168
lacosamide 200 mg twice daily | -168
more alert and responsive | -168
follow simple commands | -168
use a writing pad | -168
delirium with agitation and delusions | 0
transfer to senior behavioral health | 0
confused | 0
frail elderly female | 0
alert and oriented to self | 0
alert and oriented to month | 0
alert and oriented to year | 0
alert and oriented to location | 0
remote memory fair | 0
recent history poor | 0
perseverated on delusional beliefs | 0
leukocytosis | 0
abundant immature neutrophils | 0
empiric antibiotic treatment | 0
hyperactive delirium with agitation | 0
hypoactive delirium with significant lethargy | 24
quetiapine | 24
haloperidol | 24
risperidone | 24
mirtazapine | 48
memantine | 72
cognitive enhancer | 72
maximum daily dose | 120
minimal benefits | 120
blood cultures | 168
cerebrospinal fluid analysis | 168
meningitis/encephalitis panel | 168
paraneoplastic antibody testing | 168
cryptococcal antigen testing | 168
HIV and syphilis antibody screens | 168
urinalysis | 168
resolution of sepsis | 168
repeat EEG evaluation | 168
generalized background slowing | 168
no epileptogenic abnormalities | 168
persistent delirium | 2160
extensive nursing support | 2160
transferring | 2160
toileting | 2160
feeding herself | 2160
alert and oriented to herself | 2160
location | 2160
year | 2160
short conversations | 2160
perseverating on a particular topic | 2160
minimally interactive | 2160
poor responsiveness | 2160
discharged to long term care | 2160