28 years old | 0
female | 0
hypothyroidism | 0
hypertension | 0
polycystic ovarian syndrome | 0
presented | 0
fever | -504
myalgias | -504
nausea | -504
vomiting | -504
worked as a paramedic | 0
involved in the care of SARS-CoV-2-positive patient | -504
SARS-CoV-2 virus not detected | 0
febrile with temperature up to 105 °F | 0
upgraded to ICU | 0
palpable liver below costal margin | 0
no rash | 0
no mucosal ulcers | 0
no lymphadenopathy | 0
negative blood cultures | 0
negative urine cultures | 0
negative hepatitis B virus core IgM antibody | 0
negative hepatitis B virus surface antigen | 0
negative hepatitis C virus antibody | 0
negative hepatitis A IgM antibody | 0
positive Monospot testing for EBV | 0
elevated EBV IgM titers 46 U/mL | 0
EBV-PCR positive 552 IU/mL | 0
CT chest unremarkable | 0
CT abdomen hepatosplenomegaly | 0
liver measuring 25 cm | 0
repeat SARS-CoV-2 PCR positive | 0
transaminitis | 0
deteriorating transaminitis | 0
consultation with Hematology/Oncology | 0
concern for HLH | 0
elevated ferritin | 0
elevated fibrinogen | 0
elevated triglycerides | 0
suggested diagnostic liver biopsy | 0
suggested bone marrow biopsy | 0
declined diagnostic liver biopsy | 0
declined bone marrow biopsy | 0
not meeting all HLH criteria | 0
high suspicion for HLH | 0
started rituximab 375 mg/m2 | 0
transferred to tertiary care center | 0
fever ≥38.5 °C | 0
splenomegaly | 0
cytopenia | 0
hypertriglyceridemia | 0
elevated ferritin >500 ng/dL | 0
low or absent NK cells | 0
elevated CD25 | 0
EBV infection | 0
SARS-CoV-2 infection | 0
HLH | 0
immunosuppressive therapy | 0
dexamethasone | 0
etoposide | 0
cyclosporine | 0
rituximab | 0
tocilizumab | 0
ruxolitinib | 0
cytokine storm | 0
immunocompromised status | 0
concomitant infections risk | 0
interleukin-6 receptor blockade | 0
Janus family kinase inhibition | 0
fever persisted | 0
transferred | 0
