18 years old | 0
male | 0
history of nonalcoholic steatohepatitis | -672
alpha 1 antitrypsin deficiency | -672
underwent orthotopic liver transplant | -672
admitted to the hospital | 0
incarcerated inguinal hernia | -24
repaired uneventfully | -24
cytomegalovirus (CMV) viremia | -24
treated with valganciclovir | -24
discharged on maintenance immunosuppression | -24
presented with encephalopathy | -5
increasing home oxygen requirements | -5
required 4L nasal cannula | -5
encephalopathy characterized by sparse speech and disorientation | -5
nonfocal neurologic examination | -5
vital signs and physical examination were within normal limits | -5
white blood cell count was 9.3 × 10^9/L | -5
creatinine 2.12 mg/dL | -5
blood urea nitrogen of 53 mg/dL | -5
synthetic liver function international normalized ratio, alanine aminotransferase, aspartate aminotransferase, and bilirubin were within normal limits | -5
arterial ammonia was unusually elevated at 204 µmol/L | -5
induction dosing of intravenous ganciclovir | -5
started on empiric antibiotic coverage with vancomycin, meropenem, micafungin | -5
intravenous micronutrient supplementation for B1, B6, and levocarnitine | -5
lumbar puncture on admission revealed an opening pressure of 8 cmH2O | -5
Gram stain revealed encapsulated yeast suspicious for Cryptococcus | -5
started on liposomal amphotericin B and flucytosine | -5
started on continuous renal replacement therapy (CRRT) and rifaximin, zinc, and lactulose | -5
ammonia proceeded to unexpectedly climb to 692 µmol/L | -1
concomitant neurological deterioration necessitating mechanical ventilation | -1
empiric intravenous doxycycline | -1
urine and bronchial aspirate was obtained for Mycoplasma and Ureaplasma polymerase chain reaction (PCR) | -1
48 hours after antifungal induction and CRRT, ammonia levels had fallen to <100 µmol/L | 24
repeat lumbar punctures revealed opening pressures greater than 45 cmH2O | 24
persistent thrombocytopenia | 24
permanent CSF diversion was not possible | 24
mental status transiently improved | 24
unable to wean from mechanical ventilation | 24
require tracheostomy | 24
persistent hydrocephalus, oliguric renal failure, and progressive splenic infarcts with necrosis | 24
splenectomy | 24
magnetic resonance imaging of the brain did not reveal cytotoxic edema | 24
sepsis, duodenal leak, persisting renal failure, and failure to thrive | 24
moved to comfort care in hospice | 24
urea cycle disorder screening studies | 24
low urine orotic level | 24
normal serum citrulline and arginine level | 24