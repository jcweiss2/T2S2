37 years old | 0
primigravida | 0
twin gestation | 0
admitted to the hospital | 0
epigastric discomfort | 0
abdominal pain | 0
malaise | 0
vomiting | 0
hypertension | -168
prescribed alpha methyldopa | -168
heart rate 102/min | 0
blood pressure 170/90 mm Hg | 0
icterus | 0
foetal heart sounds heard | 0
ultra sonography of abdomen showed fatty liver | 0
ultra sonography of abdomen showed twin pregnancy | 0
haemoglobin 10.7 g% | 0
total count 10,700/mm3 | 0
platelets 2.6 lakhs | 0
urea 11 mg/dl | 0
creatinine 1.4 mg/dl | 0
uric acid 5.3 mg/dl | 0
lactate dehydrogenase 442 U/L | 0
peripheral smear negative for haemolysis | 0
hepatitis B surface antigen negative | 0
hepatitis C virus negative | 0
human immunodeficiency virus negative | 0
prothrombin time test 48 s | 0
International Normalised Ratio 4.0 | 0
total bilirubin 7.8 mg/dl | 0
direct bilirubin 4.0 mg/dl | 0
serum glutamic oxaloacetic transaminase 316 U/L | 0
serum glutamic-pyruvic transaminase 313 U/L | 0
alkaline phosphatase 974 | 0
total protein 5.3 U/L | 0
albumin 2.8 U/L | 0
globulin 2.5 U/L | 0
plasma ammonia 93 meq/d | 0
urine albumin++ | 0
cardiotocography showed evidence of foetal distress | 0
presumptive diagnosis of pre-eclampsia | 0
presumptive diagnosis of acute fatty liver of pregnancy | 0
emergency caesarean section | 0
given vitamin K | 0
given fresh frozen plasma | 0
induction by rapid sequence using thiopentone | 0
induction by suxamethonium | 0
trachea intubated | 0
anaesthesia maintained with oxygen | 0
anaesthesia maintained with Nitrous oxide | 0
anaesthesia maintained with sevoflurane | 0
anaesthesia maintained with fentanyl | 0
anaesthesia maintained with atracurium | 0
mannitol transfused | 0
albumin transfused | 0
twin babies delivered | 0
twin babies healthy | 0
extubation | 24
recovery uneventful | 24
cryoprecipitate transfused | 24
FFP transfused | 24
broad spectrum antibiotics started | 24
magnesium sulphate continued | 24
serum magnesium levels monitored | 24
liver function deteriorated | 48
tonic clonic convulsions | 72
respiratory distress | 72
mechanical ventilation initiated | 72
antibiotic changed to tobramycin | 72
computed tomography scan brain | 72
electroencephalography | 72
repeat ultra sound scan of abdomen | 72
ascites with hyperechoic features | 72
haemorrhagic ascites | 72
coagulopathy | 72
central venous pressure maintained | 72
weaned off | 168
non-invasive ventilation continued | 168
hepatic function improved | 168
viral markers negative | 168
coagulopathy corrected | 168
patient improved | 480
shifted out from post-operative intensive care unit | 480