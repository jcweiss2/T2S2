70 years old | 0
    woman | 0
    Streptococcus pneumoniae aortic valve endocarditis | -8760
    bioprosthetic porcine aortic valve replacement | -8760
    recurrent S. pneumoniae endocarditis | -8760
    aortic root replacement | -8760
    homograft | -8760
    rivaroxaban | -8760
    atrial fibrillation | -8760
    pseudomonal bacteremia | -672
    cefepime | -672
    outpatient levofloxacin | -672
    worsening right-sided chest pain | -336
    growing pulsatile mass | -336
    computed tomography angiogram | -336
    2.5 × 2.0-cm proximal thoracic aortic pseudoaneurysm | -336
    anterior mediastinal hematoma | -336
    labetalol | 0
    esmolol | 0
    prothrombin complex concentrate | 0
    vancomycin | 0
    levofloxacin | 0
    CTA 7 hours later | 7
    growth of the pseudoaneurysm to 3.4 × 2.1 cm | 7
    neck 0.6 cm wide | 7
    location 1.4 cm superior to the right coronary artery ostium | 7
    lesion was thought to be infectious | 0
    two prior sternotomies | -8760
    substernal pulsatile mass | -336
    endovascular stent graft placement | 0
    transvenous pacer | 0
    right femoral access | 0
    left axillary artery accessed | 0
    infraclavicular incision | 0
    axillary artery punctured | 0
    0.035 Glidewire | 0
    8F sheath | 0
    GLIDECATH | 0
    double-curved Lunderquist wire | 0
    pigtail catheter | 0
    left femoral 5F sheath | 0
    36 × 50-mm Zenith abdominal extension stent graft | 0
    rapid pacing | 0
    device deployed | 0
    angiography demonstrated continued pseudoaneurysm filling | 0
    stent graft angled along the lesser curve of the aorta | 0
    another 36 × 50-mm Zenith stent | 0
    completion angiography | 0
    patency of both coronary arteries | 0
    exclusion of the pseudoaneurysm | 0
    transferred to the critical care unit | 0
    antibiotic therapy changed to tobramycin | 0
    meropenem | 0
    admission blood cultures grew Pseudomonas aeruginosa | 0
    aspirin | 0
    prophylactic subcutaneous heparin | 0
    rivaroxaban discontinued | 0
    heart rate controlled with metoprolol | 0
    predischarge computed tomography scan | 240
    discharged | 240
    home infusions | 240
    2 weeks of tobramycin | 240
    6 weeks of meropenem | 240
    peripherally inserted central catheter | 240
    lifelong suppressive therapy with oral levofloxacin | 240
    follow-up CTAs at 4 months | 2880
    follow-up CTAs at 6 months | 4320
    exclusion of the pseudoaneurysm | 2880
    decreased size of the mediastinal hematoma | 2880
    stable positioning of the stent grafts | 2880
    resolution of all symptoms | 2880
    no evidence of endoleak | 2880
    infected pseudoaneurysm located at the homograft to transverse aortic arch anastomosis | -8760
    infected pseudoaneurysms often enlarge rapidly and rupture | 0
    nonoperative management likely fatal | 0
    incidence of infected aneurysms | 0
    estimates ranged from 0.7% to 2.6% | 0
    infected pseudoaneurysms treated with open surgery | 0
    endovascular intervention performed successfully | 0
    low mortality | 0
    need for reintervention | 0
    most common complications | 0
    sepsis | 0
    reinfection | 0
    Pseudomonas is a rare cause of arterial infection | 0
    high risk of the implanted stent graft to become infected | 0
    lifelong suppressive antibiotic therapy | 240
    developing endovascular solutions | 0
    short landing zones | 0
    high shear stress | 0
    left ventricular outflow tract forces | 0
    curvature of the aorta | 0
    proximity to the coronary artery ostia and arch vessels | 0
    hybrid debranching TEVAR | 0
    endovascular coiling | 0
    endovascular coiling or plugging would likely have failed | 0
    embolize the high-flow pseudoaneurysm | 0
    patient and device selection | 0
    avoid complications such as stroke and myocardial infarction | 0
    anatomic criteria for ascending aorta interventions | 0
    sinotubular junction diameter of ≤38 mm | 0
    proximal landing zone of ≥10 mm | 0
    no endovascular devices dedicated to the ascending aorta approved | 0
    studies reported successful procedures using thoracic and abdominal aortic cuffs | 0
    early data with ascending aortic devices from trials are promising | 0
    grafts from W.L. Gore & Associates | 0
    Cook Medical Inc | 0
    Bolton Medical | 0
    groups have used thoracic cuffs | 0
    advantage of easier fitting to the curvature of the aortic arch | 0
    ability to use femoral access | 0
    only used when the ascending aorta has an adequate length | 0
    limited length of the ascending aorta | 0
    14 mm of clearance above the ostia of the right coronary artery | 0
    chosen an abdominal cuff | 0
    completely covered stent | 0
    no bare metal component | 0
    length of the delivery system | 0
    ease of deployment | 0
    left axillary access | 0
    groups have favored a transapical or transcarotid approach | 0
    avoided increased stroke risk associated with transcarotid access | 0
    risk of cardiac or valvular complications with transapical approaches | 0
    graft diameter was oversized | 0
    rapid ventricular pacing | 0
    limit cardiac output and motion at the landing zone | 0
    extra care to avoid covering the coronary arteries | 0
    conversion to an open procedure likely fatal | 0
    first device landed more distally than intended | 0
    failed to exclude the pseudoaneurysm | 0
    position of the first device became advantageous | 0
    provided a scaffold to push the second device | 0
    exclusion of the pseudoaneurysm without coverage of the coronary ostia | 0
    AA-TEVAR using overlapping abdominal extension grafts | 0
    evidence that AA-TEVAR can be performed successfully | 0
    good short-term results | 0
    longer follow-up needed | 0
    durability | 0
    complications of such repairs | 0
    developing guidelines for patient and device selection | 0
    future development of devices for AA-TEVAR | 0
    branched grafts to extend the seal | 0
    devices that can be unsheathed and resheathed | 0
    aid in precise deployment | 0
    patients with a short proximal landing zone | 0
    AA-TEVAR can be performed using a second stent graft | 0
    help correctly angle another stent graft | 0
    without covering the coronary arteries | 0
    