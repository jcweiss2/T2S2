56 years old | 0
female | 0
admitted to the hospital | -1440
history of schizophrenia | -1440
perforated diverticulitis | -1440
sigmoid resection | -1440
anastomotic leak | -720
defunctioning ileostomy | -720
feculent peritonitis | -720
surgical wound dehiscence | -720
percutaneous drainage | -720
laparotomy | -720
prolonged broad-spectrum antibiotic treatment | -720
wound debridements | -720
high-protein/caloric diet | -720
acetaminophen 650 mg 4 times per day | -720
increased acetaminophen dose to 650 mg every 4 hours | -504
hypovolemic shock | 0
high gastrointestinal losses | 0
poor oral intake | 0
new abdominal collections | 0
acute kidney injury (AKI) | 0
high-anion-gap metabolic acidosis (HAGMA) | 0
elevated anion gap | 0
negative alcohol screen | 0
normal liver function tests | 0
normal lactate | 0
negative for salicylates | 0
mildly elevated beta-hydroxybutyrate | 0
elevated serum osmolal gap | 0
stopped acetaminophen | 0
started volume expansion with dextrose and bicarbonate drip | 0
N-acetyl cysteine administration | 0
sustained low-efficiency dialysis (SLED) | 0
urine organic acid testing | 24
increased excretion of 5-oxoproline | 24
improved HAGMA | 48
discharged from ICU | 48
required vasopressor and ventilatory support | 48
septic shock | 48
ventilator-associated pneumonia | 48
transferred back to the medical ward | 72
recurrent aspirations | 120
respiratory failure | 180
died | 180