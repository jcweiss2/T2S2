29 years old | 0
male | 0
cardiogenic shock | -720
biventricular failure | -720
ejection fraction 5-10% | -720
myopericarditis | -720
constrictive physiology | -720
PICC line placed | -720
discharged on milrinone | -720
fever | -24
chills | -24
septic shock | 0
PICC line removed | 0
IV vancomycin | 0
piperacillin/tazobactam | 0
vasopressor support | 0
Chryseobacterium indologenes | 48
ciprofloxacin | 48
piperacillin/tazobactam | 48
weaned off vasopressor support | 72
pericardiectomy | 216
completed 14 days of antibiotics | 336
discharged from the hospital | 360
inotrope independent | 360
follow-up | 7440
no evidence of recurrent infection | 7440
NYHA Class I | 7440
non-ischaemic cardiomyopathy | -720
viral myopericarditis | -720
constrictive pericarditis | -720
atrial flutter | -720
radiofrequency ablation | -720
inotrope therapy | -720
home milrinone infusion | -720
peripherally inserted central catheter | -720
elective pericardiectomy | -24
fever of 38.7°C | -24
tachycardia | -24
hypotension | 0
elevated lactate level | 0
blood cultures drawn | 0
Gram-negative rods | 48
infectious disease team consulted | 48
susceptibility testing | 72
sensitivity to ciprofloxacin | 72
sensitivity to piperacillin | 72
sensitivity to trimethoprim/sulfamethoxazole | 72
resistance to meropenem | 72
improved clinically | 120
afebrile | 120
negative blood cultures | 120
interval echocardiogram | 168
left ventricular EF increased | 168
right ventricular systolic dysfunction improved | 168
guideline-directed medical therapy | 360
furosemide | 360
metoprolol succinate | 360
sacubitril-valsartan | 360