70 years old | 0
male | 0
previously healthy | 0
sudden and severe loss of vision in both eyes | -96
eye pain | -96
conjunctival injection | -96
swelling | -96
oral diclofenac consumption | -144
viral prodrome | -144
rashes all over the body | -144
oral mucosal ulcerations | -144
macular rash over upper torso | 0
new ulcerating lesions over buccal and perioral tissue | 0
TEN diagnosis | 0
supportive treatment initiation in septic ICU | 0
extreme conjunctival congestion | 0
corneal sloughing | 0
corneal thinning | 0
severe anterior chamber reaction | 0
hypopyon | 0
amniotic membrane transplant planned | 0
topical moxifloxacin started | 0
lubricants started | 0
corneal perforation | 24
uveal prolapse | 24
mild proptosis | 24
lid edema | 24
restricted extraocular muscles | 24
systemic steroids | 24
electrolytes | 24
antibiotics | 24
panophthalmitis progression | 24
evisceration in both eyes | 24
death due to multi-organ failure | 72
eviscerated material sent for microbiological examination | 72
blood culture sent for microbiological examination | 72
no bacterial growth in eviscerated material | 72
no bacterial growth in blood culture | 72
