42 years old | 0
Caucasian | 0
male | 0
bilateral lung transplant | -43800
cystic fibrosis | -43800
transferred to ICU | 0
fever | 0
flu-like symptoms | 0
acute hypoxemic respiratory failure | 0
PaO2/FiO2 ratio = 81 | 0
high-flow oxygen therapy | 0
computed tomogram of the chest showed diffuse bilateral ground-glass nodular opacities | 0
areas of mosaic attenuation | 0
clinical condition deteriorated | 24
mechanical ventilation | 24
low tidal volume | 24
positive end-expiratory pressure | 24
septic shock | 24
refractory hypoxemia | 24
neuromuscular blockade with cisatracurium | 24
pulmonary vasodilator therapy with inhaled epoprostenol | 24
vasopressor support | 24
immunosuppression curtailed | 24
broad-spectrum antimicrobial therapy initiated | 24
vancomycin | 24
piperacillin-tazobactum | 24
azithromycin | 24
voriconazole | 24
prone position ventilation initiated | 24
manual proning initiated | 24
hypoxemia improvement from PaO2 81 mmHg to 168 mmHg | 24
bronchoscopic sampling deferred | 24
patient's daughter tested positive for Bordetella pertussis | 192
patient tested positive for Bordetella pertussis | 216
levofloxacin added | 216
transitioned to mechanically rotating bed | 216
prone position ventilation for 16 hours a day | 216
tolerated supine ventilation | 528
ventilator dyssynchrony | 528
deep sedation | 528
intermittent neuromuscular blockade | 528
tracheostomy | 648
liberated from mechanical ventilation | 1536
severe neuromuscular weakness | 1536
critical illness neuropathy/myopathy | 1536
ICU delirium | 1536
non-reactive pupils | 744
cessation of neuromuscular blockade | 744
neurological work-up | 744
MR imaging of the brain consistent with multifocal lesions | 744
left occipital lobe lesions | 744
central and peripheral enhancement suggesting septic emboli | 744
lumbar puncture | 744
MR angiography | 744
trans-esophageal echocardiogram | 744
serial blood cultures | 744
fundoscopic examination revealed bilateral visual loss | 744
optic nerve pallor | 744
concluded hypoxia-induced cerebral infarction | 744
increased intraocular pressure | 744
decreased ocular perfusion pressure | 744
optic nerve injury | 744
profound optic nerve pallor | 744
severe bilateral optic atrophy | 744
single A2B0 rejection | -43800
peak FEV1 post-transplant 3.32 liters (88% predicted) | -43800
pre-ICU FEV1 3.17 liters (85% predicted) | -43800
FEV1 1.74 liters (47% predicted) | 4392
legally blind from bilateral optic atrophy | 4392
retinal vascular attenuation | 4392
Bordetella pertussis pneumonia | 0
ischemic optic neuropathy | 744
