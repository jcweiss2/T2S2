60 years old | 0
male | 0
admitted to casualty | 0
bleeding from the oral cavity | 0
large clots in the oral cavity | 0
shock | 0
hemoglobin 6.1 g/dl | 0
coagulation profile normal | 0
fluid replacement | 0
blood transfusion | 0
stabilized | 0
carcinoma of hypopharynx | -8760
induction chemotherapy | -8760
concurrent chemoradiation | -8760
recurrence | -0
endoscopy | 0
large eccentric friable mass lesion in the hypopharynx | 0
bleeding | 0
CBS suspected | 0
angiography | 0
magnetic resonance angiography | 0
lesion encasing external carotid artery | 0
minimal luminal narrowing | 0
no dissection or pseudoaneurysm | 0
interventional radiologist consulted | 0
transfemoral supra-aortic digital subtraction angiogram | 0
active contrast extravasation | 0
embolization | 0
coil embolization | 0
no active extravasation of dye | 0
tiny stump of left external carotid artery | 0
successful embolization | 0
postembolization patient stable | 0
discharged | 24