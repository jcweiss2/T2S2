21 years old | 0
female | 0
admitted to the hospital | 0
dyspnea | -48
fever | -48
malaise | -48
blood pressure of 109/57 mmHg | 0
temperature of 38.2 °C | 0
heart rate of 118 bpm | 0
respiratory rate of 24 breaths/min | 0
oxygen saturation of 78% | 0
oxygen saturation improved to 97% | 0
chest X-ray demonstrated multifocal pneumonia | 0
treatment with ceftriaxone | 0
treatment with azithromycin | 0
axillary lymphadenopathy | 0
cervical lymphadenopathy | 0
inguinal lymphadenopathy |C:\Users\Acer\Documents\GitHub\KnowledgeGraphs\EventTimeline\example_case_2.tsv
respiratory decline | 0
endotracheal intubation | 0
mechanical ventilation | 0
CT chest | 0
CT abdomen | 0
CT pelvis | 0
bilateral lung consolidation | 0
moderate pericardial effusion | 0
HIV negative | 0
streptococcus pneumonia negative | 0
legionella negative | 0
histoplasma negative | 0
brucella negative | 0
aspergillus negative | 0
tuberculosis negative | 0
influenza negative | 0
respiratory syncytial virus negative | 0
mild elevation in mycoplasma IgM | 0
mild elevation in chlamydia antibody titer | 0
bronchoscopy | 0
bronchoalveolar lavage | 0
no mucus plugs | 0
no active bleeding | 0
no endobronchial lesions | 0
no anatomical abnormalities | 0
acute inflammatory cells | 0
transthoracic echocardiogram | 0
normal systolic function | 0
elevated LDH of 2319 unit/L | 0
cervical lymph node biopsy | 0
histopathology demonstrating necrotizing lymphadenitis | 0
karyorrhectic debris | 0
abundant histiocytes | 0
blood cultures negative | 0
sputum cultures negative | 0
urine cultures negative | 0
aggressive antibiotic therapy | 0
high dose steroids | 0
supportive care | 0
increasing pressure support | 0
IVIG administration | 0
hemoglobin decrease | 0
hemolytic work up | 0
haptogobin < 10 mg/dL | 0
schistocytes on peripheral smear | 0
thrombocytopenia | 0
platelet level of 26 K/mcL | 0
elevated partial thromboplastin time | 0
elevated prothrombin time | 0
elevated D-dimer levels | 0
fresh frozen plasma transfusion | 0
clinical deterioration | 0
laboratory deterioration | 0
expired | 0
DIC | 0
Kikuchi-Fujimoto disease | 0
multiorgan failure | 0
