6 years old | 0
    male | 0
    sudden onset abdominal pain | -1
    diffuse abdominal pain | -1
    vomited clear fluid twice | -1
    dehydrated tongue | 0
    diffuse abdominal tenderness | 0
    elevated white blood cell count (24,310/mm3) | 0
    nonspecific small bowel gas on plain radiograph | 0
    mild ileus | 0
    diffuse small bowel wall thickening on ultrasound | 0
    ascites on ultrasound | 0
    refused contrast-enhanced abdominal CT | 0
    discharged against medical advice | 0
    rushed to pediatric emergency department again | 15
    altered mentality | 15
    no response to painful stimuli | 15
    dilated pupils (5mm) | 15
    severe abdominal distension | 15
    uncheckable blood pressure | 15
    weakly palpable femoral pulse | 15
    percutaneous oxygen saturation (77%) | 15
    blood sugar level (22 mg/dL) | 15
    pretibial intraosseous cannulation | 15
    failure of intravenous catheterization | 15
    fluid and medications infused through intraosseous cannulation | 15
    shock state | 15
    arterial blood gas pH (7.15) | 15
    arterial blood gas bicarbonate (7.7 mM) | 15
    hemoglobin (10.1 g/dL) | 15
    hematocrit (27.7%) | 15
    rapid decrease in hemoglobin (4.7 g/dL) | 16
    rapid decrease in hematocrit (13%) | 16
    disseminated intravascular coagulopathy | 16
    antithrombin III (38.9%) | 16
    D-dimer (9.18 mg/L) | 16
    prothrombin time (1.61 INR) | 16
    activated partial thromboplastin time (43.9 seconds) | 16
    lactic acid (10.9 mmol/L) | 16
    initial hydration | 16
    central venous catheter placement via left subclavian vein | 16
    massive fluid administration | 16
    transfusions | 16
    inotropics administration | 16
    contrast-enhanced abdominal CT scan performed | 16
    systolic blood pressure maintained (90 mmHg) | 16
    large amount of ascites on CT | 16
    bowel wall thickening on CT | 16
    poor or absent enhancement of strangulated bowel segment on CT | 16
    serrated beak sign on CT | 16
    whirl sign on CT | 16
    closed loop obstruction on CT | 16
    surgical exploration | 16
    three quarters of small bowel herniated through mesenteric defect | 16
    mesenteric defect near ileocecal valve (two fingerbreadth size) | 16
    diffusely hemorrhagic small bowel | 16
    edematous small bowel | 16
    inflammatory change in small bowel | 16
    congenital internal hernia with strangulated small bowel diagnosis | 16
    resection of gangrenous small bowel (>2 meters) | 16
    anastomosis of proximal jejunum and terminal ileum | 16
    four-day treatment in pediatric intensive care unit | 96
    moved to general ward | 96
    started soft diet on 5th day post-operation | 120
    hypertension due to renal ischemic injury | 120
    short bowel syndrome | 120
    cognitive function normal | 120
    gradually improving conditions | 120