61 years old | 0
male | 0
morbid obesity | 0
Chronic Obstructive Pulmonary Disease | 0
hypertension | 0
type 2 diabetes mellitus | 0
admitted to the hospital | 0
diffusely erythematous rash | -168
rash refractory to topical nystatin therapy | -120
topical nystatin therapy | -168
erythromycin | -72
fluconazole | -72
rash spread diffusely | -72
erythematous morbilliform papules | -72
short of breath | -12
metabolic acidosis | -12
respiratory acidosis | -12
intubated | -12
hypotensive | -12
vasopressor support with norepinephrine | -12
shock liver | -12
acute kidney failure | -12
CVVHD | -12
neutrophilic leucocytosis | -12
fever | -12
discontinued erythromycin | 0
discontinued fluconazole | 0
started on broad spectrum antibiotics | 0
vancomycin | 0
meropenem | 0
micafungin | 0
discontinued antibiotics | 12
started on methylprednisolone | 12
improvement in haemodynamics | 24
improvement in rash | 24
extubated | 24
discontinued vasopressor agents | 24
recovery of kidney function | 96
recovery of liver function | 96
maintained on oral prednisone | 96
discharged | 168