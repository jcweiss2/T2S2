14 years old | 0
female | 0
diagnosed with ALL | -672
induction chemotherapy | -672
Vincristine | -672
Daunorubicin | -672
Prednisone | -672
PEG-Asparaginase | -672
pancytopenia | -4
absolute neutrophil count of 210/mm3 | -4
acute-onset left-lower-extremity pain | 0
bilateral leg pain | 4
hip pain | 4
back pain | 4
progressive weakness of both lower extremities | 4
inability to bear weight | 4
tachycardic | 4
febrile | 4
hypotensive | 4
systolic pressures in the low 80s | 4
nonspecific swelling of the left thigh | 4
tenderness of the left thigh | 4
no skin discoloration | 4
no crepitus | 4
decreases in platelet count | 4
low fibrinogen | 4
elevated thrombin time | 4
IV fluid bolus | 4
gentamycin | 4
ceftazadime | 4
left-lower-extremity Doppler ultrasound | 4
negative deep venous thrombosis | 4
necrotizing deep-soft-tissue infection | 4
General Surgery service consulted | 4
CT scan | 4
intramuscular gas in multiple muscle compartments | 4
Clostridium perfringens | 4
blood cultures | 4
operative intervention | 8
exploration and debridement | 8
extensive longitudinal incisions | 8
intact skin, subcutaneous tissue, and superficial fascia | 8
liquefactive necrosis | 8
adductor magnus involved | 8
adductor brevis involved | 8
gracilis involved | 8
gastrocnemius involved | 8
posterior hamstrings involved | 8
debridement to apparent viable tissue | 8
large defects in muscle groups | 8
Intensive Care Unit | 8
serial washouts and further debridement | 12
Vacuum-Assisted Closure device | 96
nonviable skin and subcutaneous tissue excised | 96
no sensory or voluntary motor function below knees | 120
bilateral above-knee amputations | 120
pedicled myocutaneous flaps | 120
transferred to surgical floor | 168
wounds healed well | 168
physical therapy and rehabilitation | 720
short-interval followup of two months | 720