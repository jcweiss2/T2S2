70 years old | 0
male | 0
admitted to the hospital | 0
sudden headache | 0
deteriorating consciousness | 0
resection of a pancreatic tumor | -8760
prostatic cancer | -8760
body temperature of 36.0°C | 0
heart rate of 79/min irregular | 0
blood pressure of 123/70 mmHg | 0
oxygen saturation of 100% | 0
respiratory rate of 12/min | 0
Japan Coma Scale of III-100 | 0
Glasgow Coma Scale of E1V2M5 | 0
pupils were 2 mm/4 mm | 0
light reflex was ±/± | 0
left concomitant deviation | 0
right paresis | 0
white blood cell count (WBC) of 7800/µl | 0
C-reactive protein (CRP) of 0.23 mg/dl | 0
atrial fibrillation rhythm | 0
multiple brain infarctions | 0
no thrombus detected by transthoracic echocardiography | 0
left atrial thrombus identified by transesophageal echocardiography | 24
cardiogenic cerebral infarction | 0
intubated | 12
unfractionated heparin 15,000 U administered | 12
edaravone 30 mg × 2 administered | 12
fever of 38.5°C | 48
rapid drop of blood pressure | 52
septic shock | 52
WBC 28,300/µL | 52
hemoglobin 14.3 g/dL | 52
platelet count 25.6 × 104/µL | 52
total protein 6.2 g/dL | 52
albumin 3.4 g/dL | 52
total bilirubin 0.7 mg/dL | 52
aspartate aminotransferase 22 U/L | 52
alanine aminotransferase 16 U/L | 52
lactase dehydrogenase 194 U/L | 52
alkaline phosphatase 189 U/L | 52
creatine kinase 114 U/L | 52
blood urea nitrogen 11.0 mg/dL | 52
creatinine 0.99 mg/dL | 52
C-reactive protein 1.38 mg/dL | 52
prothrombin time 79.0% | 52
activated partial thromboplastin time 66.0 s | 52
fibrinogen 686 mg/dL | 52
S. pneumoniae detected in blood and sputum cultures | 52
slight infiltration in the lower right lung field | 52
no spleen | 52
community-acquired pneumonia by Pneumococcus | 52
OPSI | 52
ceftriaxone 2 g × 2 administered | 52
IVIG 5 g × 3 days administered | 52
fluid resuscitation | 52
0.5 γ noradrenaline administered | 52
mechanical ventilation | 52
edaravone discontinued | 52
condition improved slowly | 72
catecholamines reduced | 72
extubated | 96
free from mechanical ventilation | 96
noradrenaline discontinued | 192
unfractionated heparin switched to warfarin | 192
transferred to a different hospital for rehabilitation | 216