69 years old | 0
female | 0
admitted to the hospital | 0
labile blood pressure | 0
recurrent headaches | 0
paresthesias | 0
lightheadedness | 0
decreased hearing | 0
garbled speech | 0
word-finding difficulties | 0
episodic thoracic back pain | 0
dyspnea | 0
hypertensive emergency | 0
pulmonary edema | 0
initial troponin 0.02 ng/mL | 0
troponin peaking at 6.77 ng/mL | 0
demand ischemia | 0
patent coronary arteries | 0
ECG showed non-specific anterolateral and inferior ST changes | 0
transient left bundle branch block | 0
QT prolongation | 0
moderate concentric left ventricular hypertrophy | 0
wall motion abnormalities consistent with apical ballooning syndrome | 0
akinesis of the mid- to apical left ventricular myocardium | 0
left ventricular ejection fraction (LVEF) of 37% | 0
past medical history of hypertension | -672
anxiety | -672
former smoker | -840
quit smoking | -840
denied alcohol use | 0
denied illicit drug use | 0
consumed 1–3 glasses of wine daily | -120
quit wine | -120
mother died from “heart disease” | -1000
father died from bladder cancer | -1000
brother had a stroke | -1000
family history negative for genetic syndromes | 0
history of reversible stress-induced cardiomyopathy | -2160
labile hypertension | -2160
nonspecific neurological complaints | -2160
generalized anxiety disorder | -2160
intolerance to beta-blockers | -2160
first diagnosed with takotsubo cardiomyopathy | -2628
presented to an outside hospital with chest pain | -2628
no trigger identified | -2628
echocardiogram showed an LVEF of 20% with apical dyskinesis | -2628
coronary angiogram showed minimal non-obstructive CAD | -2628
3-month follow-up echocardiogram showed complete resolution of wall motion abnormalities | -2592
normal LVEF | -2592
second episode of cardiomyopathy | -1814
presented to another outside facility with a hypertensive emergency | -1814
pulmonary edema | -1814
LVEF was again 20% with new apical dyskinesis | -1814
hyperkinetic base | -1814
no cause found | -1814
repeat echocardiogram 1 month later was normal | -1788
without wall motion abnormalities | -1788
normal LVEF | -1788
third hospital presentation | -744
nonspecific neurological complaints | -744
uncontrolled hypertension | -744
pulmonary edema | -744
labile blood pressure | -744
echocardiogram showed an LVEF of 40% with severe basal hypokinesis | -744
preserved function of the apical myocardium | -744
suggestive of reverse takotsubo | -744
repeat angiogram was unchanged | -744
CT/CTA of the chest showed no significant vascular abnormalities | -744
irregular heterogenous lesion along the left adrenal gland | -744
24-hour urine collection showed an elevated level of epinephrine | -744
normal norepinephrine | -744
normal cortisol | -744
normal dopamine | -744
home medications included a beta-blocker | 0
losartan/hydrochlorothiazide combination | 0
self-discontinued the carvedilol | -120
intolerant of metoprolol | -120
intolerant of nebivolol | -120
blood pressure was very labile | -120
difficult to control | -120
requiring multiple medication changes | -120
admitted to our facility | 0
extensive workup | 0
evaluate the cause of neurological symptoms | 0
recurrent cardiomyopathies | 0
stroke was ruled out | 0
dedicated CT and MRI scans | 0
renal artery stenosis was considered | 0
ruled out with a renal artery duplex ultrasound | 0
CTA of the chest was performed | 0
evaluate thoracic back pain | 0
hypertensive emergency | 0
no acute findings | 0
irregular heterogeneous lesion along the left adrenal gland | 0
lab work revealed normal blood counts | 0
metabolic panel | 0
thyroid function | 0
ANA | 0
negative HIV serology | 0
drug screen | 0
plasma aldosterone was normal | 0
plasma normetanephrine level was elevated | 0
plasma metanephrine was elevated | 0
thin-slice CT of the abdomen/pelvis with contrast | 0
characterize the adrenal mass | 0
7.3×4.8×7.1 cm left adrenal mass | 0
intrinsic cystic areas | 0
layering fluid | 0
measured 38 Hounsfield units (HU) on pre-contrast imaging | 0
59 HU on portal venous imaging | 0
72 HU on delayed phase imaging | 0
admitted to the intensive care unit | 0
hypertensive emergency | 0
severe anxiety | 0
managed with a nicardipine drip | 0
IV labetalol | 0
lorazepam | 0
elevated plasma metanephrines | 0
confirming the presence of an adrenal mass | 0
started on an alpha-blocker (prazosin) | 0
in addition to the labetalol | 0
uncomplicated left laparoscopic adrenalectomy | 288
performed on hospital day 12 | 288
pathology confirmed the diagnosis of pheochromocytoma | 288
postoperatively | 288
hypotensive | 288
briefly required norepinephrine | 288
recovered well from the surgery | 288
normalization of her blood pressure | 288
resolution of neurological symptoms | 288
ECG normalization | 288
discharged on post-operative day 3 | 336
on metoprolol for her cardiomyopathy | 336
seen at 1 month | 720
reported no recurrence of symptoms | 720
anxiety had greatly improved | 720
tolerating the metoprolol well | 720
repeat serum metanephrines were normal | 720
repeat echocardiogram showed normalization of the left ventricular function | 720
no residual wall motion abnormalities | 720
ECG was unremarkable | 720
seen at 6 months | 4320
reported no recurrence of symptoms | 4320
anxiety had greatly improved | 4320
tolerating the metoprolol well | 4320
seen at 12 months | 8760
reported no recurrence of symptoms | 8760
anxiety had greatly improved | 8760
tolerating the metoprolol well | 8760