43 years old | 0
male | 0
hypertension | 0
mild lacunar infarction | 0
no remnant of weakness | 0
perindopril | 0
aspirin | 0
referred for respiratory failure | 0
community-acquired pneumonia | 0
invasive ventilatory support | 0
chest X-ray consolidation right lower zone | 0
marked leukocytosis | 0
raised C-reactive protein | 0
mild hypoalbuminemia | 0
hyperglycemia | 0
normal hepatic function | 0
normal renal function | 0
normal electrolytes | 0
negative blood cultures | 0
IV co-amoxiclav | 0
transferred to ICU | 0
vital signs deterioration | 0
septic shock | 0
triple inotropes support | 0
IV piperacillin/tazobactam | 0
extubation | 168
failed oxygenation after extubation | 168
reintubation | 168
failed extubation attempts | 168
tracheostomy | 168
chest X-ray improvement | 168
persistent respiratory failure | 168
no clinical features of myasthenia gravis | 168
anti-acetylcholine receptor antibody elevated | 168
nerve conduction study decremental responses | 168
diagnosis of myasthenia gravis | 168
IV immunoglobulin | 168
pyridostigmine | 168
prednisolone | 168
azathioprine | 168
improvement after 2 weeks | 336
tracheostomy removal | 336
discharge | 336
no thymoma on CT scan | 336
Neurology Clinic follow-up | 336
no further myasthenic crises | 336
community-acquired pneumonia (previously treated) | 0
myasthenic crisis | 0
respiratory failure | 0
myasthenia gravis | 0
