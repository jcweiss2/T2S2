33 years old | 0
female | 0
Caucasian | 0
generalized anxiety disorder | 0
admitted to the hospital | 0
right ankle pain | -48
edema | -48
fall at a wedding | -48
increased edema | -24
proximal migration of edema | -24
paresthesia | -24
denies fever | -24
denies chills | -24
denies shortness of breath | -24
denies systemic symptoms | -24
elevation exacerbated pain | -24
range of motion exacerbated pain | -24
weight-bearing exacerbated pain | -24
initial X-rays | -24
no evidence of acute osseous pathology | -24
no evidence of soft-tissue gas | -24
significant edema | 0
erythema | 0
tenderness to palpation | 0
ecchymosis | 0
compartments firm but compressible | 0
mild pain with passive stretch | 0
triphasic dorsalis pedis and posterior tibial artery pulses | 0
sensation intact but diminished | 0
motor function intact | 0
referred to the emergency department | 0
venous duplex ultrasound | 0
no evidence of deep venous thrombosis | 0
admitted to the emergency room observation unit | 0
serial compartments checks | 0
initial improvement | 0
hypotensive | 12
tachycardic | 12
emergent trip to the operating room | 12
compartment releases | 12
dual incision fasciotomy | 12
dishwater fluid | 12
weakened fascia | 12
tissue biopsy | 12
fasciotomy sites copiously irrigated | 12
wound VAC placed | 12
transferred to the surgical intensive care unit | 12
norepinephrine pressors | 12
blood cultures reported positive | 12
Gram-positive cocci | 12
broad-spectrum antibiotics started | 12
vancomycin | 12
clindamycin | 12
penicillin | 12
hemodynamically unstable | 17
addition of vasopressin | 17
necrotic right foot | 17
biopsy results revealed necrotizing fasciitis | 17
right foot amputation | 17
through tibia guillotine amputation | 17
necrotic muscle, fat, and fascia | 17
guillotine amputation through the mid-thigh | 17
postoperatively stabilized | 24
managed on ceftriaxone | 24
repeat irrigation and debridement | 48
finalized above-knee amputation | 72
ambulating with a prosthesis | 6720
final X-ray | 6720