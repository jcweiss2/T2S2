58 years old | 0
female | 0
admitted to the emergency department | 0
dyspnea | 0
bilateral flank pain | 0
pallor | 0
clamminess | 0
blood pressure 170/120 mmHg | 0
heart rate 120 beats/min | 0
body temperature 38.2°C | 0
respiration rate 30 breaths/min | 0
oxygen saturation 89% | 0
body mass index 25.1 kg/m2 | 0
height 148 cm | 0
weight 55 kg | 0
phendimetrazine tartrate for weight loss | -8760
crackles in the right lung field | 0
abdomen soft without tenderness | 0
elevated CRP | 0
elevated ESR | 0
leukocytosis | 0
normocytic anemia | 0
normal platelet count | 0
suspicious acute kidney injury | 0
suspicious liver injury | 0
mixed metabolic-respiratory acidosis | 0
elevated lactate levels | 0
bilateral diffuse infiltrations on chest radiography | 0
round mass lesion in the left paravertebral area on CT | 0
sedated | 0
intubated | 0
admitted to the intensive care unit | 0
broad-spectrum antibiotics | 0
mechanical ventilation | 0
rapid resolution of lung infiltrations | 24
high fever | 0
uncontrolled hypertension | 0
elevated troponin-I | 0
elevated creatinine kinase | 0
elevated NT-proBNP | 0
hypokinetic mid inferior and apical segments on echocardiogram | 0
reduced left ventricular ejection fraction | 0
referred to an endocrinologist | 24
elevated 24-hour urinary metanephrine | 0
elevated plasma norepinephrine | 0
elevated plasma normetanephrine | 0
elevated plasma IL-6 | 0
SDHB mutation | 0
diagnosis of functional paraganglioma | 48
initiating preoperative alpha-blockers | 48
normalized body temperature | 65
controlled blood pressure | 65
open excision of the retroperitoneal mass | 408
histological examination of the tumor | 408
immunohistochemistry for chromogranin A | 408
discontinued doxazosin | 408
no postoperative complications | 408
improved inflammatory markers | 432
improved cardiac biomarkers | 432
improved renal biomarkers | 432
improved hepatic biomarkers | 432
decreased 24-hour urinary metanephrine | 432
replaced phendimetrazine tartrate with glucagon-like peptide-1 receptor agonist | 432
follow-up abdominal CT | 9360
no evidence of recurrence or distant metastases | 9360
asymptomatic during follow-up visits | 9360