74 years old | 0
male | 0
Japanese | 0
admitted to the hospital | 0
head trauma | -24
falling on a mountain | -24
no headaches | 0
no seizures | 0
no visual disorders | 0
painful bruises on arms and legs | 0
dementia | -672
Glasgow Coma Scale 13/15 | 0
heart rate 94 beats per minute | 0
blood pressure 149/75 mmHg | 0
temperature 37.9°C | 0
abrasion wound on the head | 0
bruises on the chest and upper abdomen | 0
severe tenderness in right lower leg | 0
manual muscle testing (MMT) 4/5 of right lower leg | 0
hemoglobin 13.5 mg/dL | 0
leukocyte count 19,200 cells/μL | 0
neutrophil count 15,398 cells/μL | 0
urea 25 mmol/L | 0
creatinine 0.76 mg/dL | 0
potassium 3.8 mmol/L | 0
sodium 141 mmol/L | 0
chloride 108 mmol/L | 0
creatine kinase 20,518 IU/L | 0
C-reactive protein 13.43 mg/dL | 0
tetanus vaccine administration | 0
tazobactam/piperacillin hydrate administration | 6
plain X-ray no fractures | 0
CT scan SAH, acute subdural hematoma, hypodense lesions | 0
lung and abdominal CT scans no abnormalities | 0
MR angiography no carotid stenosis, brain aneurysm, or vasospasm | 0
brain MR imaging altered intensities in bilateral parietooccipital areas | 0
hyperintense regions on T2WI, FLAIR, DWI, and ADC | 0
spinal cord MR imaging normal | 0
ascending weakness in muscles of extremities | 48
bulbar weakness | 48
complete quadriplegia | 288
bulbar palsy | 288
weakness of respiratory muscles | 288
lower oxygen saturation | 288
respiratory intubation with mechanical ventilation | 288
deep tendon reflexes (DTR) absent | 288
sensory loss not clear | 288
intravenous immunoglobulin (IVIg) administration | 288
leukocyte count 12,700 cells/μL | 288
C-reactive protein 3.50 mg/dL | 288
creatine kinase normal | 288
no anti-GM1 nor anti-GQ1b antibodies | 288
blood and cerebrospinal fluid (CSF) cultures negative | 288
IgGs of viruses not detected in CSF | 288
CSF analysis 92 mg/dL protein and 8/mmc cell count | 288
electrophysiological analysis not performed | 288
brain MR imaging increased signals of hyperintensity | 288
extubation | 576
improved MMTs of limbs | 576
brisk DTR | 576
brain MR imaging almost complete disappearance of T2WI, FLAIR, DWI, and ADC hyperintensities | 576
discharged to rehabilitation hospital | 1320