31 years old | 0
woman | 0
systemic lupus erythematosus (SLE) | 0
stage IV lupus nephritis | 0
prior stroke | -8760
intravenous drug use | 0
cardiogenic shock | 0
mental status changes | 0
three prior mitral valve replacements | -8760
recurrent nonbacterial thrombotic endocarditis (NBTE) | -8760
aggressive immunosuppression | -8760
anticoagulation | -8760
drowsy | 0
elevated jugular venous pressure | 0
prominent v wave | 0
body temperature 36.3°C | 0
blood pressure 95/66 mm Hg | 0
heart rate 94 beats/min | 0
hemoglobin 10.3 g/dL | 0
white blood cell count 18.9 × 10^9/L | 0
platelet count 64 × 10^9/L | 0
international normalized ratio 3.6 | 0
creatinine 1.7 mg/dL | 0
drug studies positive for narcotics | 0
drug studies positive for cannabis | 0
antiphospholipid serology normal | 0
blood cultures negative | 0
initiation of intravenous antibiotics | 0
diagnosis of pneumonia | 0
consideration of infectious endocarditis | 0
advised ongoing broad-spectrum intravenous antibiotics | 0
blood cultures with extended cultures | 0
serologic studies for Coxiella | 0
serologic studies for Legionella | 0
serologic studies for Chlamydia | 0
serologic studies for Bartonella | 0
serologic studies for Brucella | 0
serologic studies for Tropheryma whipplei | 0
serologic studies for HIV | 0
serologic studies for hepatitis | 0
operative cultures for Gram staining | 0
operative cultures for anaerobic and aerobic cultures | 0
operative cultures for fungal smear and culture | 0
operative cultures for acid-fast smear | 0
operative cultures for mycobacterial culture | 0
operative cultures for pathologic examination | 0
operative cultures for 16s recombinant RNA testing | 0
no culprit organisms identified | 0
transthoracic echocardiography (TTE) showing dehisced mitral valve prosthesis | 0
displaced to mid atrium | 0
severe mitral regurgitation | 0
intervalvular fibrosa completely dehisced | 0
associated cavity | 0
two dominant jets of periprosthetic regurgitation | 0
three-dimensional imaging used | 0
preoperative transesophageal echocardiography (TEE) | 0
posterior annulus dehiscence | 0
loculated cavity | 0
perivalvular regurgitation | 0
high-risk nature of planned procedure discussed | 0
decision to proceed with surgery | 0
poor clinical state | 0
young age | 0
anticipated death without intervention | 0
underwent fourth sternotomy | 0
mitral valve prosthesis dehisced along posterior annulus | 0
sitting high in left atrium | 0
close to pulmonary veins | 0
true mitral annulus displaced apically | 0
large cavity at intervalvular fibrosa | 0
multiloculations debrided | 0
surgical pathology showed bland fibrin thrombus | 0
fibrous tissue with mild chronic inflammation | 0
negative for microorganisms | 0
extensive reconstruction of fibrous skeleton of heart and atria | 0
mitral valve annulus reconstructed | 0
33-mm bioprosthesis integrated | 0
large patch of bovine pericardium used | 0
reconstruct left atrial dome | 0
reconstruct interatrial septal incision | 0
postoperative TEE showed well-seated mitral valve bioprosthesis | 0
mean gradient 3 mm Hg | 0
no regurgitation | 0
required extracorporeal membrane oxygenation | 0
left ventricular ejection fraction 25% | 0
sluggish flow in left atrium | 0
required multiple blood product transfusions | 0
postoperative day 5 TEE showed layered thrombus in left atrium | 120
underwent surgical clot removal | 120
thrombus reaccumulated in operating room | 120
extracorporeal membrane oxygenation support withdrawn | 120
patient died | 120
autopsy declined | 120
