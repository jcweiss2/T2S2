35 years old | 0
housewife | 0
gravid 3 | 0
para 2 | 0
no history of smoking | 0
no medical illness | 0
no specific medications | 0
no congenital anomalies | 0
admitted to radiology department | -28 weeks * 24 * 7 = -4704
omphalocele | -28 weeks * 24 * 7 = -4704
fetal chest with loss of anterior chest wall | -23 weeks * 24 * 7 = -3864
cardiac anomalies | -23 weeks * 24 * 7 = -3864
Pentalogy of Cantrell | -23 weeks * 24 * 7 = -3864
ectopia cordis | -23 weeks * 24 * 7 = -3864
amniocentesis not performed | -23 weeks * 24 * 7 = -3864
magnetic resonance imaging (MRI) | -23 weeks * 24 * 7 = -3864
extra-thoracic heart | -23 weeks * 24 * 7 = -3864
herniation of the left lung | -23 weeks * 24 * 7 = -3864
herniated liver | -23 weeks * 24 * 7 = -3864
dilated bowel | -23 weeks * 24 * 7 = -3864
spinal deformity | -23 weeks * 24 * 7 = -3864
parents informed | -23 weeks * 24 * 7 = -3864
ultrasonography | -33 weeks * 24 * 7 = -5544
male gender | -35 weeks * 24 * 7 = -5880
Pentalogy of Cantrell confirmed | -35 weeks * 24 * 7 = -5880
ectopia cordis confirmed | -35 weeks * 24 * 7 = -5880
caesarian section | 0
newborn length 46 cm | 0
newborn weight 2100 g | 0
head circumference 30 cm | 0
thoracic perimeter 25 cm | 0
Apgar score 3/10 | 0
Apgar score 6/10 | 5
bulky omphalocele | 0
liver and bowel loops out of the abdomen | 0
maldevelopment of the distal part of the sternum | 0
diaphragmatic hernia | 0
heart located outside the chest | 0
abnormalities | 0
admitted to neonatal intensive care unit (NICU) | 0
mechanical ventilation | 0
progressive respiratory failure | 0
severe respiratory acidosis | 0
electrolyte imbalance | 0
deteriorated general condition | 24
died on the second day | 48
septicemia | 48
respiratory failure | 48
autopsy examination not performed | 48