58 years old | 0
    female | 0
    hypertension | 0
    diabetes mellitus | 0
    Brugada syndrome | 0
    ICD implantation in 2017 | 0
    3-day febrile illness | -72
    multiple syncopal episodes | 0
    syncopal episode in 2019 | -17544
    ventricular fibrillation | -17544
    ICD shock in 2019 | -17544
    emergency department ICD interrogation | 0
    multiple episodes of ventricular fibrillation | 0
    nonsustained ventricular fibrillation | 0
    7 episodes of ventricular fibrillation | 0
    appropriate ICD shocks | 0
    fever persisted after admission | 0
    maximum temperature of 101.7°F in first 24 hours | 24
    antipyretics use | 0
    febrile periods | 0
    additional episodes of ventricular fibrillation | 24
    shock termination | 24
    rapid nasal swab positive for SARS-CoV-2 | 0
    admission to intensive care unit | 0
    isoproterenol infusion 2 μg bolus | 0
    isoproterenol infusion 1 μg/min | 0
    aggressive fever treatment with acetaminophen | 0
    aggressive fever treatment with salsalate | 0
    persistent fever | 0
    cooling blanket use | 0
    temperature normalization | 24
    no further ventricular arrhythmias | 24
    hydroxychloroquine started on day 1 | 24
    hydroxychloroquine discontinued on day 2 | 48
    QTc prolongation to 554 ms | 48
    difficult oxygenation | 0
    declining respiratory status | 0
    non-rebreather mask use | 0
    prone positioning | 0
    initial chest radiograph unremarkable | 0
    serial radiographs showing acute respiratory distress syndrome | 0
    COVID-19-associated pneumonia | 0
    isoproterenol discontinued on day 3 | 72
    atrial tachycardia with rates 140-150 bpm | 72
    broad-spectrum antibiotics started on day 5 | 120
    concern for superimposed bacterial pneumonia | 120
    remdesivir initiated on day 6 | 144
    respiratory decline requiring intubation | 144
    progressive lymphopenia 130/μL | 0
    increased C-reactive protein 54.5 mg/dL | 0
    increased D-dimer 8474 ng/mL | 0
    increased fibrinogen >1000 mg/dL | 0
    increased ferritin 1116 ng/mL | 0
    increased procalcitonin 2.7 ng/mL | 0
    therapeutic anticoagulation with LMWH | 0
    hypercoagulable state | 0
    septic shock | 0
    initiation of multiple vasopressors | 0
    infrequent atrial tachycardia | 0
    no further ventricular arrhythmias | 0
    sedation holiday on day 18 | 432
    unarousable | 432
    CT showing intracranial hemorrhage | 432
    mass effect | 432
    irreversible neurological injury | 432
    transition to comfort care | 432
    <|eot_id|>

    58 years old | 0
    female | 0
    hypertension | 0
    diabetes mellitus | 0
    Brugada syndrome | 0
    ICD implantation in 2017 | 0
    3-day febrile illness | -72
    multiple syncopal episodes | 0
    syncopal episode in 2019 | -17544
    ventricular fibrillation | -17544
    ICD shock in 2019 | -17544
    emergency department ICD interrogation | 0
    multiple episodes of ventricular fibrillation |"0
    nonsustained ventricular fibrillation | 0
    7 episodes of ventricular fibrillation | 0
    appropriate ICD shocks | 0
    fever persisted after admission | 0
    maximum temperature of 101.7°F in first 24 hours | 24
    antipyretics use | 0
    febrile periods | 0
    additional episodes of ventricular fibrillation | 24
    shock termination | 24
    rapid nasal swab positive for SARS-CoV-2 | 0
    admission to intensive care unit | 0
    isoproterenol infusion 2 μg bolus | 0
    isoproterenol infusion 1 μg/min | 0
    aggressive fever treatment with acetaminophen | 0
    aggressive fever treatment with salsalate | 0
    persistent fever | 0
    cooling blanket use | 0
    temperature normalization | 24
    no further ventricular arrhythmias | 24
    hydroxychloroquine started on day 1 | 24
    hydroxychloroquine discontinued on day 2 | 48
    QTc prolongation to 554 ms | 48
    difficult oxygenation | 0
    declining respiratory status | 0
    non-rebreather mask use | 0
    prone positioning | 0
    initial chest radiograph unremarkable | 0
    serial radiographs showing acute respiratory distress syndrome | 0
    COVID-19-associated pneumonia | 0
    isoproterenol discontinued on day 3 | 72
    atrial tachycardia with rates 140-150 bpm | 72
    broad-spectrum antibiotics started on day 5 | 120
    concern for superimposed bacterial pneumonia | 120
    remdesivir initiated on day 6 | 144
    respiratory decline requiring intubation | 144
    progressive lymphopenia 130/μL | 0
    increased C-reactive protein 54.5 mg/dL | 0
    increased D-dimer 8474 ng/mL | 0
    increased fibrinogen >1000 mg/dL | 0
    increased ferritin 1116 ng/mL | 0
    increased procalcitonin 2.7 ng/mL | 0
    therapeutic anticoagulation with LMWH | 0
    hypercoagulable state | 0
    septic shock | 0
    initiation of multiple vasopressors | 0
    infrequent atrial tachycardia | 0
    no further ventricular arrhythmias | 0
    sedation holiday on day 18 | 432
    unarousable | 432
    CT showing intracranial hemorrhage | 432
    mass effect | 432
    irreversible neurological injury | 432
    transition to comfort care | 432