34 years old| 0  
male | 0  
admitted for evaluation of penile discharge | -1008  
blurred vision in the left eye (OS) | -1008  
left knee pain of one-week duration | -1008  
Neisseria gonorrhea isolated from penile discharge | -1008  
synovial fluid aspirate was unrevealing | -1008  
presumed reactive joint inflammation | -1008  
corneal ulcer OS | -1008  
BCVA of counting fingers (CF) at 1 foot | -1008  
corneal scrapings of the ulcer | -1008  
negative for bacteria or fungi | -1008  
slit lamp examination unremarkable OD | -1008  
BCVA of 20/20 | -1008  
normal optic discs | -1008  
normal macula | -1008  
normal retinal vessels | -1008  
normal periphery in both eyes (OU) | -1008  
intensive topical treatment with moxifloxacin and natamycin every 4 hours | -1008  
healing of the corneal ulcer | -672  
rapid progressive diminution of vision OD | -336  
BCVA 20/400 OD | -336  
BCVA 20/60 OS | -336  
inferior keratic precipitates | -336  
intense anterior chamber inflammation | -336  
1-mm hypopyon | -336  
dispersed pigment on the anterior lens capsule | -336  
posterior subcapsular cataract | -336  
4+ vitreous haze | -336  
no fundus view | -336  
B scan revealed significant vitreous opacities | -336  
flat retina | -336  
healed corneal ulcer OS | -336  
large central scarring | -336  
no epithelial defect | -336  
fundus examination OS unremarkable | -336  
serum testing negative for syphilis | -336  
serum testing negative for angiotensin converting enzyme | -336  
serum testing negative for lysozyme | -336  
serum testing negative for tuberculosis (T spot) | -336  
serum testing negative for HIV | -336  
diagnosis of infective endophthalmitis suspected | -336  
urgent vitreous biopsy | -336  
pars plana vitrectomy (PPV) OD | -336  
intraoperative fundus examination revealed dense vitreous opacification | 0  
peripheral retinitis | 0  
vasculitis | 0  
localized inferotemporal rhegmatogenous retinal detachment | 0  
retinal tear | 0  
endolaser applied to the retinal tear | 0  
air-fluid exchange | 0  
aphakic | 0  
vitreous cavity filled with perfluoropropane (C3F8) | 0  
intravitreal vancomycin (1mg) | 0  
intravitreal ceftazidime (2.25 mg) | 0  
postoperative topical ofloxacin | 0  
postoperative prednisolone acetate | 0  
admitted to infectious diseases service | 0  
systemic workup for infectious source | 0  
oral levofloxacin | 0  
oral doxycycline | 0  
repeat intravitreal vancomycin (1 mg) | 48  
repeat intravitreal ceftazidime (2.25 mg) | 48  
repeat intravitreal dexamethasone (0.4 mg) | 48  
vitreous tap positive for Staphylococcus capitis | 0  
vitreous culture positive for Staphylococcus capitis | 0  
negative for toxoplasmosis | 0  
negative for lymphoma | 0  
negative for cytomegalovirus | 0  
negative for herpes simplex virus | 0  
negative for varicella zoster virus | 0  
negative for fungal agents | 0  
blood cultures negative | 0  
transthoracic echocardiography negative for vegetations | 0  
anterior chamber reaction improved | 168  
vitreous haze continued to improve | 168  
BCVA CF OD (without aphakic correction) | 504  
minimal vitreous haze | 504  
flat retina | 504  
no retinitis | 504  
50% gas fill | 504  
placement of sulcus intraocular lens | 2688  
BCVA improved to 20/80 OD | 2688  
retina remained flat | 2688  
no vitreous cavity inflammation | 2688  
<|eot_id|>
