43 years old | 0
male | 0
smoker | 0
chest pain | 0
electrocardiogram (ECG) changes suggesting postero-lateral myocardial infarction | 0
high serum troponin levels | 0
cardiac arrest (ventricular fibrillation) | 0
failed to have a return of spontaneous circulation | 0
evaluated and accepted for resuscitation with tMCS | 0
CentriMag™ Circulatory Support System introduced through left femoral artery and right femoral vein | 0
cardiorespiratory collapse reversed by tMCS via CentriMag™ within 12 minutes | 0
coronary angiogram showed severe 3-vessel coronary artery disease | 0
stents placed in two obtuse marginal arteries | 0
rest of coronary circulation unsuitable for further intervention | 0
intra-aortic balloon pump inserted | 0
left ventricular ejection fraction 19% | 0
tMCS weaning protocol suggested satisfactory recovery after 5 days | 0
neurologically intact | 0
tMCS device explanted | 120
patient suddenly deteriorated | 128
tMCS re-established via femoral approach | 128
hemodynamic status deteriorated | 360
tMCS CentriMag™ instituted again | 360
left groin sepsis | 360
arterial cannula re-sited in left subclavian artery via tube graft | 360
venous drainage via right femoral vein | 360
sepsis cleared | 0
decided to perform LVAD implantation (bridge to transplantation) | 0
continuous flow pump | 0
LVAD treatment offered | 0
type A aortic dissection confirmed by CT aortogram | 288
intimal flap extended from ascending aorta to iliac arteries | 288
no evidence of communication between true and false lumens | 288
agreed strategy prior to surgery | 0
ascending aorta replaced with tube graft | 0
Teflon strips used for distal ascending aorta | 0
myocardial protection achieved | 0
HeartMate 3 implanted | 0
HeartMate outflow graft anastomosed to aortic interposition graft | 0
weaned off cardiopulmonary bypass | 0
patient stayed in ICU for 2 weeks | 0
on ward for 4 weeks | 168
discharged home | 672
totally independent | 2928
acute type A aortic dissection repair | 0
LVAD insertion | 0
satisfactory outcome | 0
left ventricular assist device (LVAD) implantation | 0
dilated cardiomyopathy | 0
ischemic cardiomyopathy | 0
temporary mechanical circulatory support (tMCS) | 0
venoarterial extracorporeal membrane oxygenation (VAECMO) | 0
re-cannulation after weaning from VA-ECMO | 0
concomitant cardiac procedures with LVAD implantation | 0
cardiorespiratory arrest | 0
severe cardiogenic shock | 0
vascular complications | 0
witnessed cardiac arrest | 0
no major comorbidities | 0
INTERMACS profile I | 0
orthotopic cardiac transplantation unavailable | 0
long-term MCS implantation | 0
aortic dissection repair | 0
venoarterial extracorporeal membrane oxygenation (VA-ECMO) | 0
