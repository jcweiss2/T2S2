33 years old | 0
female | 0
admitted to the hospital | 0
shortness of breath | 0
feeling ill | -168
high fever | -168
tested positive for SARS-CoV-2 | -168
elevated body mass index | -672
respiratory function compromised | 0
severe hypoxemia | 0
endotracheal intubation | 0
mechanical ventilation | 0
veno-venous extracorporeal membrane oxygenation | 0
severe acute respiratory distress syndrome | 0
hemodialysis | 96
ECMO removed | 336
successful weaning | 360
impaired liver function | 0
elevated liver parameters | 0
toxic/ischemic liver injury | 0
elevated liver enzymes | 336
SSC-CIP | 336
treatment with Ursofalk | 336
computed tomography of the abdomen | 240
no signs of parenchymal damage | 240
no signs of cholestasis | 240
magnetic resonance cholangiopancreatography | 1128
mild stenosis of the distal common bile duct | 1128
suspected stricture of prepapillary CBD | 1128
endoscopic retrograde cholangiopancreatography | 1440
rarefication of intrahepatic bile ducts | 1440
SSC-CIP confirmed | 1440
magnetic resonance imaging | 3096
progressive encapsulated intrahepatic fluid accumulation | 3096
intrahepatic abscess | 3096
elevated inflammatory parameters | 1008
renal failure | 1008
hemodialysis | 1008
liver parameters remained elevated | 1008
interdisciplinary meeting | 1008
discussion of orthotopic liver transplantation | 1008
deterioration in general health | 1008
impaired respiratory function | 1008
reduced chance of successful surgery | 1008
plan for transplantation discarded | 1008
treatment with remdesivir | 0
treatment with Convalescent Plasma Transfusion | 0
treatment with antibiotics | 0
organ failure | 3696
death | 3696