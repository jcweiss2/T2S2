38 years old | 0
    woman | 0
    nondiabetic | 0
    flank pain | -120
    fever | -120
    raised total leukocyte counts | 0
    normal creatinine | 0
    significant pyuria | 0
    Escherichia coli in urine culture | 0
    10-mm obstructive calculus in left lower ureter | 0
    ureteroscopy performed | 0
    spinal anesthesia | 0
    antibiotics administered | 0
    ureteric catheter placed | 0
    thick pus drained from left pelvicalyceal system | 0
    calculus fragmented with Lithoclast | 0
    double-J stent placed | 0
    high-grade fever | 6
    hypotension | 6
    acute respiratory distress syndrome | 6
    vasopressors started | 6
    ventilator support started | 6
    transfer to intensive care | 6
    blood parameters repeated | 0
    urine culture samples taken | 0
    blood culture samples taken | 0
    piperacillin-tazobactam started | 0
    aminoglycoside started | 0
    fluid resuscitation | 0
    dopamine needed | 0
    norepinephrine needed | 0
    ventilator support in prone position | 0
    gradual improvement over 60 hours | 60
    vasopressor support for more than 5 days | 120
    ventilator support for more than 5 days | 120
    acrocyanosis of all four limbs | 0
    normal partial thromboplastin time | 0
    normal D-dimer | 0
    normal fibrinogen levels | 0
    cardiac evaluation | 0
    vasopressors continued for 3 days | 72
    acrocyanosis progressed to peripheral gangrene | 72
    multispecialty management started | 72
    plastic surgeon involved | 72
    infection disease specialist involved | 72
    anesthetists involved | 72
    antibiotic therapy continued | 72
    conservative local debridement | 72
    secondary skin grafting | 72
    sympathetic blockade attempted | 72
    left below-elbow amputation | 25 days * 24 = 600
    right below-knee amputation | 600
    loss of all fingers and toes | 600
    hospital stay for 25 days | 600
    sepsis | 0
    Gram-negative septicemia | 0
    no disseminated intravascular coagulation | 0
    