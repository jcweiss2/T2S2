57 years old | 0
male | 0
fever | -72
lumbago | -72
sudden onset persistent right flank pain | -72
fatigue | -72
fever persisted | -72
fatigue persisted | -72
right flank pain persisted | -72
admitted to the emergency room | 0
POCUS performed | 0
EPN diagnosed | 0
transferred to the ICU | 0
abdominal CT scan performed | 0
10-year history of poorly controlled diabetes | -87600
30-year history of smoking | -262800
30-year history of drinking | -262800
recent cessation of smoking and drinking | -72
temperature of 38.8 °C | 0
heart rate of 130 bpm | 0
blood pressure of 108/74 mmHg | 0
moderate dose of continuously pumped norepinephrine (0.56 μg/kg/min) | 0
respiratory rate of 22 breaths/min | 0
heart beat fast without murmurs | 0
lungs sounded clear without crackles | 0
soft abdomen | 0
abdomen not tender | 0
severe knocking tenderness in the right flank | 0
leukocytosis (10.37 × 10^9/L) | 0
neutrophils 81% | 0
hemoglobin 11.9 g/dL | 0
thrombocytopenia (69 × 10^9/L) | 0
normal alanine aminotransferase (21 IU/L) | 0
normal aspartate aminotransferase (23 IU/L) | 0
normal bilirubin (0.58 mg/dL) | 0
elevated serum creatinine (1.66 mg/dL) | 0
increased C-reactive protein (175.1 mg/L) | 0
elevated procalcitonin (> 100 ng/mL) | 0
glycosylated hemoglobin 9% | 0
heavy pyuria (325/μL) | 0
arterial blood gas pH 7.43 | 0
partial pressure of carbon dioxide 36.8 mmHg | 0
partial pressure of oxygen 64.4 mmHg | 0
bicarbonate 24.8 mmoL/L | 0
elevated lactate level 2.9 mmoL/L | 0
positive blood culture for extended spectrum beta-lactamase-producing Escherichia coli | 0
positive urine culture for Escherichia coli | 0
emergency POCUS on day 3 showing hyperechoic foci with dirty shadowing and comet-tail artifacts | 0
"falls" sign identified | 0
abdominal CT scan confirming EPN | 0
gas collection in right perirenal space | 0
enlarged right kidney with perinephric fat stranding | 0
mild right hydronephrosis | 0
absence of urinary stones | 0
fluid resuscitation | 0
insulin infusion | 0
vasopressor support | 0
broad-spectrum antibiotic therapy (meropenem and tigecycline) | 0
repeat CT scan on day 7 showing abscess and more perinephric fat stranding | 168
CT-guided PCD performed on day 5 | 120
pus culture yielding E. coli | 120
discontinuation of norepinephrine within 5 days | 120
CT reexaminations on days 9 and 11 showing catheter placement and gas/abscess absorption | 216, 264
asymptomatic with normal serum creatinine | 216, 264
normal platelet count | 216, 264
perirenal catheter removed | 336
discharged on day 14 | 336
oral levofloxacin prescribed | 336
repeat urinary CT scan at 2 weeks post-discharge showing normal kidney imaging | 672
stable blood glucose control during follow-up | 13176
normal renal function during follow-up | 13176
patient satisfied with care | 13176
