57 years old | 0
    female | 0
    hypertension | 0
    recurrent cystitis | 0
    type 2 diabetes mellitus | 0
    ESRD on hemodialysis (3 sessions/week) | 0
    brought into the emergency room | 0
    found lethargic | -12
    barely conscious | -12
    previous hospital admissions for recurrent UTI | 0
    previous hospital admissions for bacteremia | 0
    last hemodialysis session | -48
    temperature of 95.5F | 0
    heart rate 102 beats per minute | 0
    respiratory rate 10 cycles per minute | 0
    blood pressure 76/55 mmHg | 0
    soft abdomen | 0
    mild distension | 0
    trace pedal edema | 0
    difficult to assess for rebound tenderness | 0
    intubated | 0
    admitted to the MICU | 0
    leukocytosis | 0
    normocytic anemia | 0
    lactic acidosis | 0
    elevated serum creatinine levels | 0
    hemoglobin A1C level 6.1% | 0
    arterial blood gas levels normal | 0
    urinalysis positive for bacteria | 0
    urinalysis positive for leukocyte esterase | 0
    urinalysis positive for nitrites | 0
    abdominopelvic CT scan extensive small and large bowel thickening | 0
    abdominopelvic CT scan no evidence of obstruction | 0
    abdominopelvic CT scan no evidence of perforation | 0
    thickening and irregularity of the bladder wall | 0
    mild ascites | 0
    abdominopelvic CT scan 1 year prior circumferential thickening of the bladder wall | -8760
    chest X-ray normal | 0
    brain CT scan normal | 0
    initiated on intravenous fluids | 0
    empiric IV antibiotics (Vancomycin and Tazobactam/Piperacillin) | 0
    norepinephrine for septic shock | 0
    continuous renal replacement therapy | 0
    general surgery team consulted for possible complicated ischemic colitis | 0
    surgical team presumptive diagnosis of ischemic colitis | 0
    surgical team presumptive diagnosis of bacteremia | 0
    no acute surgical intervention warranted | 0
    persistently febrile | 24
    tachycardic | 24
    requiring more doses of norepinephrine | 24
    abdomen more distended | 24
    laboratory parameters significantly worsened | 24
    blood microbiology studies resulted for Escherichia coli | 24
    urine microbiology studies resulted for Escherichia coli | 24
    taken to the operating room for exploratory laparotomy | 48
    necrotic bladder wall | 48
    ruptured bladder wall | 48
    free fluid in the abdominopelvic cavity | 48
    no bowel ischemia | 48
    no bowel perforation | 48
    partial cystectomy | 48
    pathologic analysis confirmed bladder tissue inflammation | 48
    pathologic analysis confirmed necrosis | 48
    no malignancy | 48
    family decided to withdraw life support treatment | 144
    died | 156
    