57 years old | 0
male | 0
mechanic | 0
medical history of occasional use of cocaine | 0
gradually worsening vision | -120
optic nerve atrophy | -120
tripped over a low brick wall | -1
fell about one meter on the back of his head | -1
tetraplegic | -1
transferred to a level 1 trauma center | 0
complete cord lesion on the level of C3 and C4 | 0
congenital narrowing of the spinal canal at the level of C3 and C4 | 0
old fracture of the third thoracic vertebra | 0
hemorrhage in the myelum at the level of C3 and C4 | 0
transferred to the Intensive Care Unit | 0
ventilator support | 0
acute respiratory distress syndrome (ARDS) | 72
pneumonia in the right lower lobe | 72
aspiration | 72
purulent sputum | 72
Haemo-lytic Streptococcus group C | 72
Streptococcus pneumoniae | 72
Haemophilus influenzae | 72
Enterobacter cloacae | 72
piperacillin/tazobactam | 72
percutaneous tracheostomy | 240
weaning | 240
no longer dependent on ventilator support | 480
discharged to a rehabilitation center | 1824
admitted again | 2628
fever | 2628
diarrhea | 2628
productive cough | 2628
pulmonary tuberculosis | 2628
Mycobacterium tuberculosis | 2628
tuberculostatic triple therapy | 2628
pseudomembranous colitis | 2628
Clostridium toxins | 2628
metronidazol | 2628
free of diarrhea | 2638
deep venous thrombosis | 2700
erysipelas | 2700
ulceration on the fingers | 2700
Escherichia coli | 2700
Klebsiella pneumoniae | 2700
Pseudomonas aeruginosa | 2700
Morganella morganii | 2700
Proteus mirabilis | 2700
urine positive for Klebsiella pneumoniae | 2700
urine positive for Enterococcus faecalis | 2700
surgically treated | 2700
heterozygosity in MBL2 exon 1 | 0
heterozygosity in MBL2 promoter region Y-221X | 0
homozygosity for the minor allele in MASP2 Y371D | 0
heterozygosity in FCN2 T236M | 0
heterozygosity in FCN2 A258S | 0
homozygosity for the minor allele in TLR2 T-16934A | 0
heterozygosity in CD14 C-159T | 0