39 years old | 0
male | 0
admitted to the hospital | 0
presented to the emergency department | 0
progressive epigastric pain | -168
nausea | -168
vomiting | -168
constipation | -168
rectal adenocarcinoma (13 years ago) | -113832
abdomino-perineal resection (13 years ago) | -113832
end colostomy surgery (13 years ago) | -113832
adjuvant chemoradiation therapy (13 years ago) | -113832
fever (39°C) | 0
tachycardia (145 bpm) | 0
hypotension (BP 90/50 mmHg) | 0
generalized abdominal tenderness | 0
guarding | 0
rebound tenderness | 0
leukocytosis (18,500 WBC/cm³) | 0
anemia (Hb 8.6 mg/dL) | 0
pneumoperitoneum on chest X-ray | 0
nil by mouth | 0
IV fluid resuscitation | 0
IV broad-spectrum antibiotics | 0
generalized peritonitis | 0
emergency laparotomy | 0
ileum perforation | 0
purulent fluid in peritoneal cavity | 0
ileum resection | 0
anastomosis | 0
abdominal cavity washout with saline | 0
significant adhesions | 0
hemodynamic instability | 0
transferred to ICU | 0
intubation | 0
imipenem | 0
tazocin | 0
vancomycin | 0
caspofungin | 0
continuous norepinephrine infusion | 0
fentanyl for pain | 0
sedation | 0
maintenance IV fluid therapy | 0
cardiac arrest | 36
CPR | 36
intensive fluid resuscitation | 36
clinical improvement | 36
extubation (day 5) | 120
clinical deterioration (day 7) | 168
febrile | 168
triple contrasted abdominal CT | 168
colo-splenic fistula | 168
splenectomy | 168
left hemicolectomy | 168
moderately differentiated adenocarcinoma | 168
necrosis | 168
viable adenocarcinoma in spleen | 168
return of intestinal peristalsis | 168
increased appetite | 168
resolved septic status | 168
discharged | 960
follow-up at one month | 720
follow-up at three months | 2160
follow-up at six months | 4320
annual surveillance colonoscopy | 8760
ulcerated mass in right colon | 8760
adenocarcinoma confirmed | 8760
total colectomy | 8760
end ileostomy insertion | 8760
