35 years old | 0
    male | 0
    intermittent crampy abdominal pain | -2160
    hypogastrium pain | -2160
    weight loss | -2160
    stools decreased in consistency | -2160
    abdominal ultrasound (multiple heterogeneous liver lesions, splenomegaly) | -720
    carcinoembryonic antigen elevation | -720
    CA 19-9 antigen elevation | -720
    computerized axial tomography (metastatic liver lesions, colon thickening, descending colon tumor) | -720
    admission to General Hospital of Mexico | 0
    abdominal pain (10/10) | 0
    fever | 0
    unstable vital signs | 0
    hypotension | 0
    tachycardia | 0
    respiratory distress | 0
    abdominal distension | 0
    generalized pain | 0
    involuntary muscular resistance | 0
    positive rebound | 0
    bowel sounds of metallic hue | 0
    leukocytosis | 0
    neutrophilia | 0
    anemia | 0
    thrombocytosis | 0
    hyperglycemia | 0
    uremia | 0
    creatinine elevation | 0
    hyperuricemia | 0
    hypocholesterolemia | 0
    hypertriglyceridemia | 0
    hyperbilirubinemia | 0
    elevated liver enzymes | 0
    hypoalbuminemia | 0
    hypoproteinemia | 0
    elevated lactic dehydrogenase | 0
    electrolyte abnormalities | 0
    coagulopathy | 0
    elevated procalcitonin | 0
    metabolic acidosis | 0
    elevated lactate | 0
    abdominal X-ray (intestinal dilation, inter-loop edema) | 0
    chest radiograph (subdiaphragmatic free air) | 0
    exploratory laparotomy | 0
    colonic perforation | 0
    left colon tumor | 0
    ascending colon tumor | 0
    para-aortic ganglionic chain invasion | 0
    free intestinal fluid | 0
    liver metastases | 0
    abscesses | 0
    radical total colectomy | 0
    Brooke-type terminal ileostomy | 0
    hemodynamic instability | 0
    septic shock | 0
    multiple organ failure | 0
    ileostomy functioning | 12
    refractory septic shock | 48
    cardiorespiratory arrest | 48
    death | 48
    