32 years old | 0
female | 0
ventriculoperitoneal shunt (VPS) | 0
weakness in bilateral upper and lower limbs | -336
altered sensorium | -336
pineocytoma | -4320
obstructive hydrocephalus | -4320
right frontal burr hole | -4320
endoscopic third ventriculostomy | -4320
ventriculoperitoneal shunting | -4320
radiotherapy | -720
headache | -504
vomiting | -504
generalized seizures | -48
admission to ICU | -24
difficulty in moving limbs | -24
febrile | 0
conscious | 0
Glasgow Coma Score (GCS) 4/15 | 0
diminished deep tendon reflexes | 0
CT scan brain revealed heterogeneous lesion | 0
residual tumor | 0
trans ependymal CSF seepage | 0
fasting blood sugar 126 mg/dl | 0
random blood sugar 289 mg/dl |*0
shunt tapped | 0
ventricular fluid with 20 RBC/mm³ | 0
ventricular fluid with 40 WBC/mm³ | 0
glucose 79 mg/dl | 0
protein 71.4 mg/dl | 0
gram-positive cocci on gram stain | 0
shunt externalized | 0
extraventricular device placed | 0
Staphylococcus lugdunensis resistant to penicillin | 0
susceptible to all other antibiotics tested | 0
afebrile | 72
discharged | 240
reinternalization of VPS | 240
follow-up to neurosurgery OPD | 720
