63 years old | 0
male | 0
presented to the emergency department | 0
midepigastric pain | -72
intolerance to oral intake | -72
denied hematemesis | 0
denied hematochezia | 0
denied other gastrointestinal symptoms | 0
midepigastric tenderness | 0
computed tomography scan | 0
fluid collection along the undersurface of a thickened duodenum wall | 0
infrarenal saccular abdominal aortic aneurysm | 0
no evidence of free air | 0
esophagogastroduodenoscopy | 0
abnormal mucosa | 0
possible mass | 0
perforation of the third portion of the duodenum | 0
taken to the operating room | 0
gross contamination from intestinal fluid | 0
perforation of the posterior medial aspect of the second portion of the duodenum | 0
saccular mycotic aortic aneurysm | 0
aortic wall inflammation | 0
aortic wall thinning | 0
impending rupture | 0
pancreaticoduodenectomy | 0
open abdominal aortic aneurysm repair | 0
rifampin-soaked Dacron graft | 0
omental wrap | 0
staged Whipple reconstruction | 48
pancreatic ductal adenocarcinoma | 0
extension through the duodenum wall | 0
lymph nodes positive | 0
margins uninvolved | 0
intractable intra-abdominal sepsis | 0
died | 3840