31 years old | 0  
    female | 0  
    non-smoking | 0  
    Caucasian | 0  
    no past medical history | 0  
    sudden-onset severe headache | -840  
    left arm numbness | -840  
    postpartum | -840  
    cranial computed tomography (CT) scan | -840  
    grade 2 subarachnoid hemorrhage (Hunt and Hess scale) | -840  
    no prior history of head injury | -840  
    uncomplicated pregnancy | -840  
    uncomplicated vaginal delivery | -840  
    admitted to the neurosurgical ward | -840  
    digital subtraction angiography (DSA) | -840  
    ruptured right middle cerebral artery aneurysm | -840  
    percutaneous endovascular coil embolization | -840  
    no permanent neurological deficits | -840  
    postpartum endometritis | -840  
    fever | -840  
    chills | -840  
    constant abdominal pain | -840  
    purulent uterine discharge | -840  
    denied urinary symptoms | -840  
    denied respiratory symptoms | -840  
    blood culture samples obtained | -840  
    empiric antibacterial therapy | -840  
    piperacillin/tazobactam | -840  
    vancomycin | -840  
    azithromycin | -840  
    sepsis | -840  
    septic shock | -840  
    transferred to the intensive care unit | -840  
    body temperature 38.3°C | 0  
    invasive blood pressure 90/65 mmHg | 0  
    crystalloid administration | 0  
    vasopressor administration | 0  
    heart rate 135/min | 0  
    arterial oxygen saturation 82% | 0  
    mild disorientation | 0  
    slower capillary refill | 0  
    coarse rales over lower lung zones | 0  
    SOFA score 4 | 0  
    hemoglobin 6.8 g/dL | 0  
    d-dimers 4.58 μg/mL | 0  
    C-reactive protein 322 mg/L | 0  
    fibrinogen concentration 6.4 mL | 0  
    E. coli sensitive to piperacillin/tazobactam | 0  
    chest radiography | 0  
    pulmonary nodules up to 40 mm | 0  
    CT thorax confirmation | 0  
    diagnostic work-up for gestational trophoblastic neoplasia | 0  
    transvaginal ultrasound | 0  
    enlarged uterus | 0  
    complete loss of zonal anatomy | 0  
    abdominal MRI | 0  
    enlarged heterogenous myometrial mass | 0  
    splenic metastatic lesion | 0  
    serum β-hCG 232,085 mUI/mL | 0  
    suction evacuation | 0  
    curettage | 0  
    choriocarcinoma diagnosis | 0  
    FIGO score 12 | 0  
    term pregnancy | 0  
    <4 months interval from pregnancy to chemotherapy | 0  
    β-hCG 97,521 mIU/mL | 0  
    >8 metastatic lesions | 0  
    brain metastasis (oncotic aneurysm) | 0  
    largest tumor lesion within the lung 40 mm | 0  
    chemonaïve | 0  
    metastatic choriocarcinoma | 0  
    high risk of resistance to single-drug chemotherapy | 0  
    multiagent chemotherapy regimen initiated | 0  
    low-dose etoposide 100 mg/m2 | 0  
    cisplatin 20 mg/m2 | 0  
    clinical improvement | 168  
    EMA/CO regimen | 168  
    etoposide | 168  
    methotrexate | 168  
    actinomycin D | 168  
    cyclophosphamide | 168  
    vincristine | 168  
    six cycles completed | 168  
    β-hCG levels plateaued | 168  
    restaging with MRI brain | 168  
    18F-FDG PET/CT scan | 168  
    decreased pulmonary nodules | 168  
    decreased uterine mass | 168  
    SUV <3.8 | 168  
    revised FIGO score 7 | 168  
    β-hCG 6 mIU/mL | 168  
    <4 metastatic lesions | 168  
    largest lesion <3 cm | 168  
    prior multiagent chemotherapy | 168  
    EP/EMA regimen | 168  
    etoposide plus cisplatin | 168  
    normalization of β-hCG | 168  
    free of disease for two years | 168  
    grade 3 neutropenia | 168  
    granulocyte colony stimulating factor (G-SCF) | 168  
    dose reduction of etoposide | 168  
    dose reduction of actinomycin D | 168  
    grade 2 alopecia | 168  
    grade 2 nausea | 168  
    dexamethasone | 168  
    ondansetron | 168  
    grade 2 fatigue | 168  
    use of male condoms | 168  
    chemotherapy toxicity | 168  
    treatment delays avoided | 168  
    unplanned pregnancy prevented | 168  