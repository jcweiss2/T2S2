52 years old | 0
female | 0
admitted to the hospital | 0
shortness of breath | 0
exacerbation of heart failure | 0
echocardiogram | 0
aortic root dilated ascending aorta | 0
bicuspid aortic valve | 0
moderate mixed aortic valve disease | 0
mild mitral regurgitation | 0
penicillin allergy | -672
Bentall’s procedure | -672
bio-integral valve aortic bio-conduit | -672
mitral valve annuloplasty | -672
sternal wound healed | -12
discharging sternal sinus | -48
infection of the sternal wires | -48
Staphylococcus aureus | -48
chronic sternal osteomyelitis | -48
sternal wound debridement | -48
removal of the superior infected sternal wires | -48
antibiotics | -48
negative pressure wound therapy | -48
conventional dressings | -48
co-trimoxazole | -48
chest pain | -24
dizziness | -24
active bleeding from her sternal wound | -24
hematoma | -24
anemia | -24
raised inflammatory markers | -24
CT angiogram | -24
pseudoaneurysm at the distal anastomosis of the ascending graft | -24
aorto-cutaneous fistula | -24
multidisciplinary team meeting | -24
endovascular stent graft | -24
Valiant Navion stent graft | -24
deployment of the stent graft | -24
completion angiogram | -24
CT angiogram after the procedure | 48
infectious disease team | 48
long-term antibiotics | 48
cardiothoracic clinic appointments | 336
vascular clinic appointment | 1008
repeat CT angiography | 1008
community nurse visits | 1008
dietician assessments | 1008
regular blood tests | 1008
red blood cell transfusions | 1008
iron infusions | 1008
psychological input | 1008
psychiatric input | 1008
social work input | 1008
septic shock | 2016
blood pressure | 2016
heart rate | 2016
respiratory rate | 2016
temperature | 2016
white cell count | 2016
C-reactive protein | 2016
lactate | 2016
CT angiogram | 2016
new infected pseudoaneurysm | 2016
multidisciplinary meeting | 2016
thoracic endovascular aortic repair | 2016
extension of the graft | 2016
intraoperative transesophageal echocardiogram | 2016
second ascending stent graft | 2016
deployment of the stent graft | 2016
completion angiogram | 2016
CT angiogram after the procedure | 2024
sternal wound bleeding | 2772
hemoptysis | 2772
dizziness | 2772
CT angiography | 2772
extension of the pseudoaneurysm | 2772
empyema | 2772
palliation | 2772
death | 3024