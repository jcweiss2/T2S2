50 years old | 0
unremarkable medical history | 0
admitted to the emergency department | 0
fever | -120
acute respiratory failure | 0
febrile for 5 days | -120
rapidly worsening shortness of breath | -24
dry cough | -24
chest x-ray performed in the ED | 0
bilateral multifocal involvement of the lungs | 0
marked diffuse interstitial pattern | 0
mildly elevated white blood cells | 0
increased C-reactive protein | 0
low procalcitonin | 0
denied recent travel history | 0
denied close contacts with animals | 0
denied contacts with sick people | 0
denied intravenous drugs use | 0
cigarette smoke | 0
frequent unprotected heterosexual intercourse | 0
tachypnea | 0
fever (101°F) | 0
hypotension | 0
tachycardia | 0
diminished vesicular breath sounds | 0
unremarkable physical examination | 0
suspicion of Pneumocystis jirovecii pneumonia | 0
HIV-1 antibody-antigen test positive | 0
weak positivity for pneumococcal urinary antigen | 0
severe hypoxemia | 0
high oxygen supply with reservoir bag | 0
blood cultures | 0
empirical therapy with piperacillin-tazobactam | 0
levofloxacin | 0
cotrimoxazole | 0
transferred to the intensive care unit | 0
mechanical ventilation | 0
bronchoscopy | 96
Gram stain of bronchoalveolar lavage negative | 96
no bacterial growth on BAL cultures | 96
no fungal growth on BAL cultures | 96
P jirovecii negative | 96
cotrimoxazole ceased | 96
no acid-fast bacteria | 96
Mycobacterium tuberculosis-complex PCR negative | 96
cytomegalovirus negative | 96
Epstein-Barr virus negative | 96
herpes simplex virus 1/2 negative | 96
adenovirus negative | 96
influenza A/B nucleic acid amplification negative | 96
Aspergillus galactomannan antigen negative | 96
BAL cytology: macrophages 32% | 96
neutrophils 63% | 96
lymphocytes 5% | 96
no neoplastic cells | 96
pneumococcal urinary antigen test repeated | 96
pneumococcal urinary antigen test negative | 96
blood cultures negative | 96
Legionella urinary antigen negative | 96
serology for intracellular bacteria negative | 96
repeated bronchoscopy | 144
Gram stain negative | 144
Ziehl-Neelsen stain negative | 144
no bacterial growth on BAL cultures | 144
no fungal growth on BAL cultures | 144
Pneumocystis jirovecii IFA negative | 144
PCR-mediated tests for viruses negative | 144
procalcitonin repeated twice | 144
procalcitonin 0.5-0.6 ng/mL | 144
no clinical improvement | 168
no radiological improvement | 168
persistently febrile | 168
severe respiratory distress | 168
control chest x-rays persistently showed interstitial bilateral pattern | 168
acute respiratory distress syndrome radiological signs | 168
confirmatory HIV Western blot negative | 24
HIV Western blot repeated | 120
Fiebig stage IV | 120
plasma HIV-RNA >10000000 cps/mL | 120
CD4+ T-cell count 571 cells/mm3 | 120
CD8+ T-cell count 234 cells/mm3 | 120
CD4+/CD8+ ratio 2.44 | 120
previous negative HIV test 6 months before admission | -4320
HIV-RNA on BAL 206647 cps/mL | 192
ART introduced | 192
tenofovir disoproxil fumarate/emtricitabine | 192
darunavir/ritonavir 800/100 mg | 192
raltegravir 400 mg bid | 192
worsening respiratory failure | 192
septic shock | 192
noradrenaline | 192
neutrophilia | 192
increased CRP | 192
chest x-ray unchanged | 192
bronchoaspirate positive for KPC-Kp | 192
high-dose meropenem | 216
gentamicin | 216
tygeclicine | 216
blood cultures negative | 216
hemodynamically stable | 216
progressive improvement of respiratory distress | 216
control chest x-rays showed improvement | 336
extubated | 336
transferred to the pneumology ward | 336
transferred to the infectious diseases unit | 432
oxygen supply de-escalated | 432
clinical improvement | 432
follow-up bronchoscopy | 648
BAL cultures positive for KPC-Kp | 648
HIV-RNA on BAL 177 cps/mL | 648
ART well tolerated | 648
discharged | 816
plasma HIV-RNA 97 cps/mL | 1344
plasma HIV-RNA <40 cps/mL | 2016
