29 years old | 0 | 0 
female | 0 | 0 
admitted to the hospital | 0 | 0 
complex regional pain syndrome | -8760 | 0 
sports-related injury | -8760 | -8760 
shoulder surgery | -8760 | -8760 
recurrent shoulder infections | -8760 | -120 
Pseudomonas aeruginosa | -8760 | -120 
Sphingomonas paucimobilis | -8760 | -120 
Candida colliculosa | -8760 | -120 
Staphylococcus aureus | -8760 | -120 
left shoulder tendon release and revision | -720 | -720 
development of CRPS | -720 | 0 
severe pain | -720 | 0 
allodynia | -720 | 0 
edema | -720 | 0 
muscle spasms | -720 | 0 
temperature changes | -720 | 0 
electromyography evaluation | -120 | -120 
brachial plexus injury | -120 | -120 
asthma | -8760 | 0 
selective IgG3 deficiency | -8760 | 0 
oral medical management | -120 | 0 
opioids | -120 | 0 
antidepressants | -120 | 0 
antispasmodics | -120 | 0 
left stellate ganglion blockade | -168 | -168 
continuous cervical epidural infusions | -168 | -168 
decreased pain | -168 | -168 
improved participation with physical therapy | -168 | -168 
reduction in oral opioid requirements | -168 | -168 
placement of a left C6–C7 interlaminar epidural catheter | 0 | 0 
fluoroscopic guidance | 0 | 0 
preprocedure labs | 0 | 0 
complete blood count | 0 | 0 
complete metabolic panel | 0 | 0 
creatinine phosphokinase | 0 | 0 
antibiotic prophylaxis | -1 | 0 
vancomycin | -1 | 0 
intrathecal and intravascular placement | 0 | 0 
lidocaine | 0 | 0 
epinephrine | 0 | 0 
epidural infusion | 0 | 120 
bupivacaine | 0 | 120 
hydromorphone | 0 | 120 
clonidine | 0 | 120 
oral home medications | 0 | 120 
methadone | 0 | 120 
diazepam | 0 | 120 
baclofen | 0 | 120 
amitriptyline | 0 | 120 
decrease in pain | 0 | 24 
less muscle spasms | 0 | 24 
increased infusion | 24 | 24 
demand dose | 24 | 120 
improved sleep | 24 | 120 
further decrease in LUE spasms and edema | 24 | 120 
febrile | 120 | 120 
wean the infusion | 120 | 120 
remove the epidural catheter | 120 | 120 
progressive headache | 120 | 120 
neck pain | 120 | 120 
increase in temperature | 120 | 120 
neurological examination | 120 | 120 
blood and urine cultures | 120 | 120 
chest x-ray | 120 | 120 
laboratory workup | 120 | 120 
increase in white count | 120 | 120 
cephalosporin | 120 | 120 
cefepime | 120 | 120 
abatement of fever | 120 | 120 
decrease in white count | 120 | 120 
MRI of the cervical spine | 120 | 120 
epidural collection | 120 | 120 
compression of the left C5 and C6 nerve roots | 120 | 120 
effacement of the thecal sac | 120 | 120 
interstitial edema in the left paraspinal muscles | 120 | 120 
transfer to the neurosciences intensive care unit | 120 | 120 
hourly neurological examination | 120 | 144 
intractable nausea and vomiting | 144 | 144 
left arm weakness | 144 | 144 
emergent decompression and evacuation | 144 | 144 
C3 to C7 cervical laminectomies | 144 | 144 
C4–C5 and C5–C6 left foraminotomies | 144 | 144 
intraoperative cultures | 144 | 144 
P aeruginosa | 144 | 144 
susceptible to cefepime | 144 | 144 
vancomycin stopped | 144 | 144 
cefepime continued | 144 | 144 
resolution of arm weakness | 144 | 216 
uneventful postoperative course | 144 | 216 
discharged home | 216 | 216 
intravenous cefepime | 216 | 1008