85 years old | 0
female | 0
admitted to the hospital | 0
painful swelling | 0
bilateral submandibular | 0
submental | 0
upper neck areas | 0
edematous skin | 0
reddish skin | 0
ill-defined reddish border | 0
extreme pain | 0
fever | 0
body temperature of 39 | 0
endodontic treatment | -72
odontogenic abscess | 0
steroid treatment | -672
arthralgia | -672
WBC of 10.26×10^3/µL | 0
ESR of 3 mm/hr | 0
neutrophil of 93.1% | 0
aPTT of 45.9 seconds | 0
CRP of 202.96 mg/L | 0
CT scan | 0
disseminated deep neck abscess | 0
left submandibular space | 0
upper mediastinum | 0
anterior neck space | 0
supraclavicular area | 0
axillary area | 0
incision and drainage | 0
necrotic fascia | 0
fasciitis | 0
triple antibiotic regimen | 0
penicillin | 0
aminoglycoside | 0
metronidazole | 0
silicon drains | 0
microscopic examination | 0
acute and chronic infection | 0
lymphocyte infiltrations | 0
necrotic fascia | 0
pus culture | 0
betahemolytic streptococcal infection | 0
sensitive to most antibiotics | 0
condition not improved | 96
CT scan | 96
infection spread | 96
under the trapezius muscle | 96
intense hot and reddish skin | 96
airway obstruction | 96
WBC of 13.18×10^3/µL | 96
ESR of 15 mm/hr | 96
neutrophil of 87.7% | 96
aPTT of 46.3 seconds | 96
CRP of 151.46 mg/L | 96
drainage under the trapezius muscle | 96
tracheostomy | 96
artificial airway | 96
ventilator therapy | 96
skin infection extended | 240
upper chest | 240
shoulder area | 240
follow-up CT images | 240
multifocal abscess | 240
left chest wall | 240
carotid area | 240
WBC of 12.21×10^3/µL | 240
ESR of 11 mm/hr | 240
neutrophil of 75.7% | 240
aPTT of 38.6 seconds | 240
CRP of 14.2 mg/L | 240
uncontrolled NF | 240
third operation | 240
incision on the chest | 240
necrotic tissue | 240
fasciotomy | 240
vancomycin monotherapy | 240
Actinibacter baumanni | 240
resistant to cabepenem | 240
infection decreased | 288
skin necrosis | 288
distal clavicular area | 288
bilobed rotational flap | 888
tracheostomy tube removed | 960
discharged | 1056
WBC of 10.08×10^3/µL | 1056
ESR of 5 mm/hr | 1056
neutrophil of 71.3% | 1056
aPTT of 25.7 seconds | 1056
CRP of 20.4 mg/L | 1056