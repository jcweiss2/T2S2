66-year-old|0
man|0
dual-chamber pacemaker implanted|0
sick sinus syndrome|0
paroxysmal atrial fibrillation|0
severe lumbar back pain|0
deteriorated rapidly|0
mental status changes|0
hypotension|0
acute renal failure|0
hypoxemic respiratory failure|0
emergent intubation|0
severe sepsis|0
hemodynamic support with vasopressin|0
hemodynamic support with norepinephrine|0
blood cultures yielded methicillin-sensitive Staphylococcus aureus|0
empirically started on vancomycin|0
antibiotic coverage narrowed to nafcillin|0
transthoracic echocardiogram demonstrated left ventricular ejection fraction of 55%|0
positive bubble study|0
patent foramen ovale|0
Doppler demonstrated medium-sized patent foramen ovale measuring approximately 2.99 cm|0
computed tomography scan revealed osteomyelitis of the lower spine (L2–L3)|0
magnetic resonance imaging demonstrated multiple small acute infarctions|0
septic emboli to the distal extremities|0
repeat blood cultures revealed the same organism for 3 consecutive days|0
transesophageal echocardiogram (TEE) performed|0
long (0.26 × 3.6 cm) mobile structure within the right atrium|0
vegetation|0
second mobile structure attached to the pacemaker lead within the right ventricle|0
no evidence of aortic and/or mitral valve endocarditis|0
no evidence of aortic arch infected atheromata|0
consulted cardiothoracic surgery|0
deemed a poor surgical candidate|0
hemodynamic instability|0
decision to perform laser lead extraction|0
concerns about septic pulmonary embolism|0
fragmentation of the vegetation leading to further cerebral and systemic emboli|0
devised system to debulk/remove vegetations|0
arrived in the hybrid operating room|0
intubated and sedated|0
bilateral femoral veins accessed|0
16F GORE® DrySeal Flex introducer sheath placed in the right common femoral vein|0
8F sheath inserted into the left common femoral vein|0
9F sheath placed in the right femoral vein|0
8F catheter (CARTO SoundStar) advanced into the right atrium|0
12F 45-degree curved sheath advanced into the right atrium|0
115-cm Indigo CAT8 XTORQ advanced into the right atrium|0
intracardiac echocardiography (ICE) used|0
vegetation attached to the RV lead with the stalk at the tricuspid valve level|0
aspiration performed with vacuum pump generating -20 inHg|0
two aspiration passes with 100 mL drawn each|0
intraprocedural ICE revealed no lingering vegetation|0
strained blood revealed presence of smaller vegetation|0
second pass performed|0
strained blood revealed large vegetation|0
Indigo Penumbra system withdrawn into the inferior vena cava|0
laser lead extraction performed|0
RA and RV leads successfully extracted|0
pocket inspected and closed with suture|0
Penumbra and ICE systems removed|0
hemostasis achieved|0
procedure time 72 minutes|0
blood loss 200 mL|0
vegetations sent to pathology|0
gram staining showed gram-positive cocci in chains|0
culture-positive for methicillin-sensitive Staphylococcus aureus|0
patient's condition improved for the first 48 hours|48
patient's condition deteriorated after 72 hours|72
tissue necrosis of the distal upper and lower extremities|72
lactic acidosis|72
worsening renal failure|72
family decided to withdraw care|72
patient extubated to comfort care|72
patient died|72
