54 years old | 0
male | 0
frontotemporal dementia | -120 months
apathy | -120 months
self-destructive impulsivity | -120 months
bedridden | - months 
weakness of lower limb | - months
frequent syncope | - months
fluctuation of blood pressure | - months
anticholinergic drug | - months
severe atrophy of bilateral frontal and temporal lobes | - months
selective serotonin reuptake inhibitors | - months
anticonvulsants | - months
dopamine agonist | - months
anticholinergic medications | - months
anemia | 0
bleeding of stomach cancer | 0
hemoglobin 8.3 g/dl | 0
atrial fibrillation | 0
admitted to the hospital | 0
subtotal gastrectomy | 0
thiopental 170 mg | 0
vecuronium 6 mg | 0
intubated | 0
mechanical ventilation | 0
sevoflurane | 0
stable vital signs | 0
systolic/diastolic BP 110–130/70–90 mmHg | 0
HR 80–95 beats/min | 0
sudden drop in BP to 70/40 mmHg | 2
shedding 300 ml of blood | 2
atrial fibrillation at varying rates between 110–130 beats/min | 2
volume of 1,500 ml of Lactated Ringer's solution | 2
1 unit of packed red blood cells | 2
TEE | 2
normal valves and contractility with adequate volume state | 2
no regional wall motion abnormality | 2
estimated ejection fraction was 65% | 2
synchronized cardioversion at 50 J | 2
HR returned to 50 beats/min | 2
no change in BP | 2
bolus injection of ephedrine | 2
infused dopamine of 10 µg/kg/min | 2
infused dobutamine of 10 µg/kg/min | 2
infused norepinephrine of 0.3 µg/kg/min | 2
no response to those drugs | 2
high dose of epinephrine at 0.5–1.0 mg | 2
increasing BP | 2
vasopressin at a rate of 4 units/h | 2
bolus dose of 10 units | 2
BP and HR returned to baseline values | 2
BP 110/65 mmHg | 2
HR 75 beats/min | 2
dopamine of 5 µg/kg/min | 2
dobutamine of 5 µg/kg/min | 2
arginine vasopressin at a rate of 4 U/h | 2
operation completed successfully | 4
transferred to the intensive care unit | 4
all vasopressors were titrated | 24
stopped completely | 24
extubated | 24
transferred to the general ward | 48
no sequelae | 48