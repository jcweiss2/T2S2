101 years old | 0
male | 0
admitted to the hospital | 0
cough | -24
productive sputum | -24
wheezing | -24
hypertension | 0
coronary artery disease | 0
old cerebral infarction | 0
diabetes mellitus | 0
no recent travel to populated areas | 0
stayed at home for months | 0
WBC 9.28×10^9/L | 0
neutrophils 80.4% | 0
lymphocytes 11.3% | 0
C-reactive protein (CRP) 2.67 mg/dl | 0
Procalcitonin (PCT) <0.05 ng/mL | 0
CT scan of the lung showed new patchy ground glass opacities | 0
community acquired pneumonia | 0
received regular infection treatment with flomoxef and levofloxacin | 0
fever | 48
adenovirus IgM positive | 48
meropenem and tigecycline prescribed | 48
no significant improvement in body temperature | 504
clinical condition began to deteriorate | 504
persistent fever | 504
lethargy | 504
thrombocytopenia | 504
elevated creatinine and transaminase levels | 504
remarkable increase in PCT | 504
antibiotic treatment switched to vancomycin and piperacillin/tazobactam | 504
respiratory failure | 864
CT scan of the chest revealed new bilateral patchy infiltrates | 864
lung cavity (7 mm × 8 mm) in the anterior segment of the left upper lobe | 864
bronchoscopy performed | 864
yellowish-white secretion almost blocked the lumen of the left main bronchus | 864
mucosa was edematous and congested | 864
samples collected from the anterior segment of the left upper lobe by bronchoalveolar lavage | 864
mNGS analysis of the BALF revealed the presence of E. faecium | 888
E. faecium with 10, 376 sequences | 888
pathogen identification confirmed by BALF culture | 888
isolate found to be resistant to vancomycin | 888
isolate sensitive to linezolid | 888
linezolid (600 mg IV q12d) started | 888
clinical condition improved | 936
platelets dropped sharply | 936
linezolid discontinued | 1008
contezolid (400 mg PO q12d) started | 1008
thrombopoietin administered | 1008
clinical improvement noted | 1056
platelet counts returned to normal | 1056
cavitary lesion resolved | 1056
patchy infiltrations decreased | 1056
contezolid therapy continued for nearly 4 months | 1056
contezolid well tolerated | 1056
platelet levels remained relatively stable | 1056
follow-up CT scan performed | 2304
lung cavity lesion and patchy infiltrations completely disappeared | 2304
contezolid discontinued | 2304