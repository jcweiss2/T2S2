42 years old | 0
female | 0
brought in due to sudden onset altered mental status | 0
low grade fevers | -120
sudden deterioration in mental status | 0
history of intravenous drug use | -10560
extraction of all maxillary teeth | -3240
mandibular dental infection | -2160
oral amoxicillin | -2160
temperature 36.7 °C | 0
heart rate 98 beats/min | 0
respiratory rate 17 breaths/min | 0
blood pressure 131/66 mm Hg | 0
oxygen saturation 99% | 0
denied fevers | 0
denied chills | 0
denied chest pain | 0
denied dyspnea | 0
denied nausea | 0
denied vomiting | 0
denied diarrhea | 0
denied skin lesions | 0
denied numbness | 0
denied tingling | 0
denied weakness of the lower extremities |8|0
holosystolic murmur at the apex | 0
petechial rash scattered on the abdomen | 0
petechial rash on palms | 0
petechial rash on soles of the feet | 0
encephalopathy | 0
facial droop | 0
slurred speech | 0
admitted to intensive care unit | 0
empiric antibiotic treatment with vancomycin | 0
empiric antibiotic treatment with meropenem | 0
unresponsive to voice | 24
minimally responsive to pain | 24
left hemi-neglect | 24
right gaze deviation | 24
Glasgow Coma Scale 6 | 24
intubated for airway protection | 24
leukocytosis 24.7 × 109/L | 0
87.6% neutrophils | 0
platelet count 17 × 109/L | 0
normal liver function | 0
normal kidney function | 0
declined HIV test | 0
acute to subacute embolic infarcts in cerebral hemispheres | 0
acute to subacute embolic infarcts in cerebellar hemispheres | 0
largest infarct involving right lentiform nucleus | 0
largest infarct involving corona radiata | 0
proximal right internal carotid artery T-shaped acute thrombus | 0
occlusion of the right middle cerebral artery | 0
subarachnoid hemorrhage in right parietal region | 0
subarachnoid hemorrhage around posterior aspect of midbrain | 0
echo densities on tricuspid valve | 0
echo densities on aortic valve | 0
echo densities on mitral valve | 0
valvular vegetations | 0
blood culture grew S. marcescens | 0
S. marcescens pansensitive susceptible to ceftriaxone | 0
S. marcescens susceptible to cefepime | 0
S. marcescens susceptible to ceftazidime | 0
S. marcescens susceptible to meropenem | 0
S. marcescens susceptible to gentamicin | 0
S. marcescens susceptible to tobramycin | 0
S. marcescens susceptible to amikacin | 0
S. marcescens susceptible to ciprofloxacin | 0
S. marcescens susceptible to levofloxacin | 0
antibiotic changed to cefepime | 72
cardiothoracic surgery consulted | 72
poor candidate for surgery | 72
neurological status deterioration | 144
no cough reflex | 144
no gag reflex | 144
fixed pupils | 144
mid-dilated pupils | 144
withdrawal of care | 144
discharged to hospice care | 144
triple valves involvement | 0
innumerable emboli | 0
severe neurological sequelae | 0
diagnosed with infective endocarditis | 0
septic embolization to the brain | 0
numerous infarcts | 0
sub-arachnoid hemorrhage | 0
denied weakness of the lower extremities | 0
leukocytosis 24.7 × 10^9/L | 0
platelet count 17 × 10^9/L | 0
