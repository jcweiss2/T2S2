21 years old | 0
male | 0
admitted to the hospital | 0
shortness of breath | -120
fever | -120
sore throat | -120
empiric treatment with vancomycin | 0
empiric treatment with piperacillin-tazobactam | 0
empiric treatment with azithromycin | 0
endotracheal intubation | 0
hypoxemic respiratory failure | 0
acute respiratory distress syndrome (ARDS) | 0
bilateral pulmonary infiltrates | 0
thrombophlebitis of the left internal jugular vein | 0
blood cultures grew Fusobacterium necrophorum | 0
blood cultures grew Granulicatella | 0
septic thrombophlebitis (Lemierre syndrome) | 0
antibiotics narrowed to piperacillin-tazobactam | 72
vancomycin restarted | 72
repeated sampling of the respiratory system for cultures | 72
sputum culture on hospital day 1 identified normal respiratory flora | 24
BAL specimens on hospital days 3 and 7 revealed no growth | 72
febrile with persistent leukocytosis | 120
empyemas with bilateral pneumothoraces | 168
surgical chest tube insertions | 168
bacterial culture performed on pleural fluid demonstrated growth of Mycoplasma hominis | 168
azithromycin therapy restarted | 168
fevers subsided | 216
liberated from mechanical ventilation | 408
discharged from the hospital | 504
Fusobacterium taxa identified by 16S rRNA gene sequencing | 0
Mycoplasma taxa identified by 16S rRNA gene sequencing | 0
whole metagenome sequencing (WMGS) performed | 0
Mycoplasma hominis identified by WMGS | 0
Fusobacterium necrophorum identified by WMGS | 0
plasma biomarkers measured | 0
RAGE measured | 0
IL-6 measured | 0
procalcitonin measured | 0
NGS data analyzed | 0
antibiotic management decisions made | 0