28 years old | 0
male | 0
farmer | 0
ingestion of two fresh tablets of Celphos | -4
vomiting | -4
abdominal pain | -4
agitated | 0
anxious | 0
irritable | 0
pulse rate not palpable | 0
blood pressure not recordable | 0
heart rate 110/min | 0
respiratory rate 28/min | 0
oxygen saturation 95% | 0
sinus tachycardia | 0
T wave inversion in lead 3 | 0
intravenous crystalloids | 0
IV magnesium sulphate | 0
IV calcium gluconate | 0
IV hydrocortisone | 0
IV dopamine | 0
noradrenaline | 0
gastric lavage with potassium permanganate | 0
activated charcoal | 0
metabolic acidosis | 0
pH 7.2 | 0
HCO3 8 mmol/L | 0
PCO2 33 mmol/L | 0
intubated | 0
shifted to ICU | 0
blood pressure 60-80 mmHg | 6
pulse rate 120/min | 6
respiratory rate 20/min | 6
input/output 3L/300 ml | 24
monomorphic ventricular tachycardia | 48
DC cardio-version | 48
IV amiodarone | 48
cardiac bio-markers raised | 48
normal sinus rhythm | 48
pH 7.4 | 96
HCO3 18 mmol/L | 96
CO2 42 mmol/L | 96
blood urea 100 mg/dl | 96
serum creatinine 4.5 mg/dl | 96
urine output 400 ml/24 hours | 96
AST/ALT 80/90 IU/L | 96
ALP 200 U/L | 96
S bilirubin 2.5 mg/dl | 96
liver and kidney involvement | 96
blood pressure 100/70 mmHg | 120
pulse rate 110/min | 120
respiratory rate 22/min | 120
total leucocyte count 14000/mm3 | 120
polymorphonuclear leucocytosis | 120
urea 200 mg/dl | 120
S. creatinine 7.5 mg/dl | 120
urine output 400 ml/24 hours | 120
pH 7.1 | 120
HCO3 10 mmol/L | 120
haemodialysis | 120
haemodialysis | 168
blood urea 70 mg/dl | 168
creatinine 4.0 mg/dl | 168
urine output 1200 ml/24 hours | 168
extubated | 144
shifted to step down unit | 192
vitals normal | 192
liver and kidney functions improving | 192
discharged | 336