84 years old | 0
female | 0
admitted to the hospital | 0
chronic kidney disease | 0
hypertension | 0
mild cognitive dysfunction | 0
uterine mass | 0
fever | -48
dry cough | -48
dyspnea | -48
heavy rain | -48
bilateral lower lung patches | 0
pleural effusion | 0
septic shock | 0
acute kidney injury | 0
respiratory failure | 0
antibiotics | 0
fluid resuscitation | 0
tracheal intubation | 0
transferred to a tertiary hospital | 0
admitted to the intensive care unit | 0
curved gram-negative bacteria isolated from blood culture | 0
direct gram stain of the pleural fluid demonstrated curved gram-negative bacilli | 0
oxidase-positive | 0
catalase-negative | 0
urease-negative | 0
glucose-nonfermenting | 0
VITEK MS failed to identify the bacterium | 0
VITEK2 GN ID card reported Burkhoderia mallei with 90% probability | 0
diagnosis of infection caused by Paludibacterium species | 0
16S rRNA polymerase chain reaction (PCR) assay | 0
primers 11F and 1512R used to amplify the conserved 16s rRNA genes | 0
1.5-kb amplified fragments from blood and pleural effusion cultures identified as Paludibacterium purpuratum | 0
pleural effusion culture did not yield any bacteria | 0
16S rRNA sequencing for the inoculated broth identified the existence of P. purpuratum | 0
pneumonia and empyema responded well to ampicillin-sulbactam | 0
bilateral pleural drainage with 24-Fr chest tubes | 0
extubated | 96
acute kidney injury resolved | 96
discharged home | 480
analyses of 16S rRNA gene sequences showed that the clinical P. purpuratum blood isolate shared the highest sequence similarity with P. purpuratum KJ031 | 0
whole-genome sequencing of the P. purpuratum strain B53371 | 0
genome size for the P. purpuratum strain B53371 is 3.63 M | 0
morphology, drug susceptibility, and metabolic abilities were assayed for the P. purpuratum B53371 strain | 0
P. purpuratum isolate was able to grow on blood agar plate and chocolate agar plates at 35°C | 0
gram stain showed curved and long gram-negative bacilli | 0
indole test for P. purpuratum isolate was negative | 0
hanging drop motility test showed a negative result | 0
isolate grew less at 42°C than that at 35°C | 0
did not grow on MacConkey plate or colistin nalidixic acid blood agar plate | 0
colony morphology on blood agar plate was small and gray at 24 hours | 0
colony morphology on blood agar plate became smooth, translucent, or white at 48 hours | 0
colony morphology on chocolate agar plate showed a white or translucent appearance at 48 hours | 0
isolated strain showed low minimal inhibitory concentration (MIC) levels for ampicillin/sulbactam, piperacillin/tazobactam, cefotaxime, cefepime, fluoroquinolones, meropenem, and aminoglycosides | 0
high MIC level for colistin in vitro | 0
phenotype microarray plates were used to analyze the metabolic profiles of the P. purpuratum strain | 0
strain was able to ferment carbon, nitrogen, phosphorus, and sulfur substrates | 0
test strain could utilize 33 substrates, mainly carbon- and nitrogen-containing sources | 0
infection might have acquired through inhalation of pathogens stirred by heavy rainfall | 0
P. purpuratum could be misidentified by the VITEK2 GN ID card diagnostic system | 0
probability for Burkholderia mallei was only 90% | 0
P. purpuratum and B. mallei share similar morphology features on blood agar and chocolate plates | 0
cultivation of this facultatively anaerobic Paludibacterium is susceptible to an array of antibiotics in vitro except for colistin | 0
whole-genome sequencing analysis revealed that the P. purpuratum isolate carried ICR-Mo, a chromosomally encoded determinant of colistin resistance | 0
ICR-Mo encodes an enzyme that helps to modify lipid A by transferring phosphoethanolamine moiety from its donor phosphatidylethanolamine to the 1’- (or 4’)-phosphate position of lipid A | 0
expression of ICR-Mo in bacteria may prevent the formation of reactive oxygen species induced by colistin | 0
present case recovered well with ampicillin/sulbactam therapy | 0
first invasive P. purpuratum infection in Taiwan | 0
infection in susceptible hosts might happen due to exposure or inhalation of this pathogen accidentally | 0