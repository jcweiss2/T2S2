67 years old | 0\
female | 0\
body weight 50 kg | 0\
height 158 cm | 0\
admitted to the hospital | 0\
backache | -672\
calculi in both kidneys associated with ureteral calculi | -672\
HLL combined with double J catheterization | -672\
purulent urine | -672\
fever | -0.5\
chill | -0.5\
low blood pressure | -0.5\
imipenem and Cilastatin sodium | -0.5\
fluid resuscitation | -0.5\
Norepinephrine | -0.5\
Hydrocortisone sodium succinate hormone | -0.5\
anuric | -48\
ARDS | -48\
invasive ventilatory support with endotracheal intubation | -48\
CRRT | -48\
transferred to the ICU | -48\
sedated state | 0\
blood pressure 80/62 mmHg | 0\
Norepinephrine 1.5 μg/kg/min | 0\
Epinephrine 1.0 μg/kg/min | 0\
heart rate 139 beats/min | 0\
transcutaneous oxygen saturation 80% | 0\
cold, clammy extremities | 0\
loud bubbling sound in the lung | 0\
oxygen partial pressure 50 mmHg | 0\
lactic acid 10.6 mmol/L | 0\
bicarbonate 10.8 mmol/L | 0\
central venous pressure 20 cmH2O | 0\
B lines in the lung | 0\
diffuse dysfunction | 0\
LVEF 20.3% | 0\
sinus tachycardia | 0\
broad ST depression | 0\
troponin I 10.2 ng/mL | 0\
amino-terminal brain natriuretic peptide precursor >35,000 pg/L | 0\
creatinine 356 μmol/L | 0\
anuria | 0\
VA-ECMO treatment | 0\
ECMO venous leading-out end used a 20F catheter | 0\
arterial leading-in end used a 17F catheter | 0\
No. 6 arterial catheter was placed in the right femoral artery | 0\
ECMO ran normally 3000 rpm | 0\
blood flow 3.5 L/min | 0\
arterial pressure 135 mmHg | 0\
venous pressure −29 mmHg | 0\
Norepinephrine stopped | 0.5\
Epinephrine stopped | 0.5\
CRRT | 0.5\
Imipenem and Cilastatin sodium combined with Vancomycin | 0.5\
lactic acid level declined | 2\
vasoactive drugs completely stopped | 10\
arterial blood lactate level normal | 12\
extended-spectrum β-lactamase-positive Escherichia coli | 48\
inflammatory indices diminished | 48\
anti-infection regimen continued | 48\
minimum serum trough concentration of Vancomycin 15–20 μg/mL | 48\
LVEF 35% | 120\
black and necrotic skin | 120\
successfully weaned from ECMO therapy | 144\
renal function scaled as acute kidney injury grade 3 | 144\
bedside CRRT discontinued | 144\
urinating | 144\
vascular ultrasonography and computed tomography angiography | 168\
vascular surgery consultation | 168\
necrotic tissues of the lower extremity amputated | 336\
spontaneous breathing successful | 120\
trachea opened | 240\
anti-infective therapy replaced by Cefoperazone sodium and Sulbactam sodium | 240\
bedside physical rehabilitation started | 240\
weaned from the ventilator | 480\
tracheotomy tube sealed | 600\
discharged | 768\
intermittent hemodialysis | 768\
take care of herself | 2160\
intermittent hemodialysis | 2160