25 years old | 0
female | 0
head-on motor vehicle collision | -1
located in the center rear passenger seat | -1
single transverse band seat belt | -1
hemodynamically stable | 0
patent airway | 0
Glasgow Coma Scale of 15 | 0
Focused Abdominal Sonography for Trauma (FAST) scan | 0
perisplenic fluid | 0
pelvic fluid | 0
no solid organ injury | 0
no pneumoperitoneum | 0
lower left rib fractures | 0
compression fractures | 0
anterior wedging of L1 and L2 | 0
transverse process fracture | 0
conservative management | 0
admitted to the Intensive Care Unit (ICU) | 0
acutely hemodynamically unstable | 72
physical examination findings concerning for an acute abdomen | 72
repeat FAST scans showing increase in free intraperitoneal fluid | 72
septic shock | 72
exploration | 72
retroperitoneal hematoma | 72
steatonecrosis plaques | 72
incomplete jejunal laceration | 72
complete section of the pancreas | 72
peripancreatic hematoma | 72
necrohemorrhagic pancreatitis | 72
distal pancreatectomy | 72
splenectomy | 72
jejunal enterorraphy | 72
open abdomen | 72
open abdomen management | 72
catastrophic abdomen | 120
complex enterocutaneous fistulas | 120
aspiration probes | 120
Goretex mesh | 120
linitud films | 120
short-gut syndrome | 2160
home parenteral nutrition | 2160
discharged | 2592
abdominal reconstruction | 8760
elective surgery | 8760
re-establish the intestinal transit | 8760
en bloc excision | 8760
subtotal colectomy | 8760
resection of the intestinal ileostomy | 8760
excision of three segments of the small intestine | 8760
reconstruction of the intestinal transit | 8760
permacol mesh plasty | 8760
wide skin flap | 8760
discharged | 8784
follow-up control | 10512
without incidents | 10512