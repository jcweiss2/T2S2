69 years old | 0
    male | 0
    hyperlipidemia | 0
    hypertension | 0
    bioprosthetic mitral valve replacement | -8760
    left parietal hemorrhage | -336
    left middle cerebral artery stroke | -336
    thrombectomy | -336
    sedation | -336
    intubation | -336
    external ventricular drain placement | -336
    mild fatigue | -336
    headache | -336
    warfarin | 0
    aspirin | 0
    rosuvastatin | 0
    holosystolic murmur III/IV at apex | 0
    no peripheral stigmata of endocarditis | 0
    mobile echodensities on posterior mitral valve leaflet | 0
    cefepime (2g IV every 8 hours) | 0
    gentamicin (80mg IV every 8 hours) | 0
    vancomycin (1250mg IV twice daily) | 0
    Aspergillus galactomannan antigen elevation | 0
    1,3-β-D-glucan elevation | 0
    Aspergillus fumigatus detected by Karius test | 0
    liposomal amphotericin B (3mg/kg IV every 24 hours) | 0
    voriconazole (360mg PO twice daily) | 0
    Aspergillus fumigatus culture positive | 144
    fungal endophthalmitis (right eye) | 144
    intravitreal voriconazole (100mcg) | 144
    valve repair surgery deferred | 144
    switch to isavuconazole (372mg daily) | 504
    therapeutic isavuconazole levels | 504
    discharge to inpatient rehabilitation | 792
    switch to micafungin (150mg IV daily) | 1200
    renal insufficiency (creatinine increase 0.34mg/dL) | 1200
    worsening generalized weakness | 1920
    failure to thrive | 1920
    elevated white blood cell count (14.3 K/UL) | 1920
    splenic infarcts | 1920
    splenic abscess | 1920
    renal infarcts | 1920
    vancomycin added (1250mg IV) | 1920
    cefepime added (2g IV every 8 hours) | 1920
    hypotension requiring vasopressors | 1944
    persistent mobile echodensity on mitral valve | 1944
    elevated 1,3@-β-D-glucan | 1944
    elevated galactomannan antigen | 1944
    acute embolic occlusions in lower extremities | 1944
    thrombectomy | 1944
    worsening hypoxemia requiring intubation | 1944
    mechanical ventilation | 1944
    increased vasopressor requirements | 1944
    transition to comfort measures | 1944
    death | 1944