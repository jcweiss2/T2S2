10 years old | 0
male | 0
admitted to the hospital | 0
kidney transplantation | -168
end-stage kidney disease | -168
PU valves | -120
vesico-ureteric reflux | -120
resection of PU valves | -72
bilateral ureteric reimplantation | -72
growth retardation | -168
underweight | -168
mother donated kidney | -168
induction therapy | -168
triple immunosuppression | -168
tacrolimus | -168
prednisolone | -168
mycophenolate sodium | -168
prophylaxis for pneumocystis | -168
prophylaxis for cytomegalovirus | -168
high fever | -48
severe cough | -48
vomiting | -48
no loss of smell | -48
no loss of taste | -48
no diarrhea | -48
normal urine output | -48
weight 22.5 kg | 0
temperature 101°F | 0
respiration 26/min | 0
pulse 120/min | 0
blood pressure 120/80 mm Hg | 0
SpO2 92% | 0
throat normal | 0
chest clear | 0
graft kidney nontender | 0
rapid antigen test positive | 0
nasopharyngeal swab sent | 0
HRCT chest CORADS-6 | 0
TSS 18/25 | 0
normal urinalysis | 0
Hb 11.3 g/dL | 0
lymphocytes 820 cells/mm3 | 0
serum creatinine 0.5 mg/dL | 0
SGPT 48 U/L | 0
CRP 9.3 mg/L | 0
ferritin 203 ng/mL | 0
LDH 403 U/L | 0
procalcitonin 0.11 ng/mL | 0
D-dimer 201 ng/mL | 0
ultrasound scan normal | 0
doppler study normal | 0
blood cultures sent | 0
throat swabs sent | 0
tacrolimus trough levels analyzed | 0
qt-PCR for CMV analyzed | 0
qt-PCR for BK virus analyzed | 0
adequate hydration | 0
antipyretics | 0
piperacillin-tazobactam | 0
RT-PCR for SARS-CoV-2 positive | 24
tacrolimus continued | 24
prednisolone continued | 24
mycophenolate stopped | 24
remdesivir administered | 24
afebrile | 144
mild cough | 144
oxygen saturations normal | 144
urine output normal | 144
creatinine stable | 144
liver functions normal | 144
PCR for CMV negative | 144
PCR for BK virus negative | 144
blood cultures sterile | 144
throat swab cultures sterile | 144
discharged | 192
home-quarantine | 192
telehealth follow-up | 192
asymptomatic | 360
renal functions normal | 360
lymphocyte count normal | 360
CRP normal | 360
HRCT chest TSS 3/25 | 360
mycophenolate restarted | 360