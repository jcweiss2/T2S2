49 years old | 0
male | 0
admitted to the hospital | 0
cough | -504
fever | -504
emaciation | -504
mass on the left side of the neck | -168
mass below the right side of the chin | -168
treated with ceftazidime | -168
fever resolved | -168
mass on the neck grew | -168
physical examination | 0
body temperature of 38°C | 0
two palpable masses | 0
inflamed and sensitive to touch | 0
moist rales in the upper lobe of the left lung | 0
white blood cell count of 14,200 cells/µL | 0
neutrophil count of 12,200 cells/µL | 0
lymphocyte count of 1.39 cells/µL | 0
platelet count of 167,000/µL | 0
hemoglobin of 124 g/L | 0
C-reactive protein level of 167.04 mg/L | 0
erythrocyte sedimentation rate of 70 mm/h | 0
procalcitonin of 0.61 ng/mL | 0
total CD3+, CD4+, and CD8+ T-lymphocyte counts | 0
liver and kidney function test results were normal | 0
level of total immunoglobulin was within the normal limit | 0
galactomannan index was 0.35 | 0
HIV negative | 0
CT of the neck revealed mixed-density lesions | 0
started on ceftazidime and levofloxacin | 0
resection of the neck masses | 24
pus sample was sent for culture | 24
B. cepacia was cultured from the mass on the neck and submental pus | 168
drug sensitivity test | 168
continued administration of ceftazidime and levofloxacin | 168
fever resolved | 168
masses decreased in size | 168
productive cough | 336
CT showed that the neck masses shrank | 336
exudative consolidation shadow in the left upper lobe | 336
left hilar lymphadenopathy | 336
bronchofibroscopy revealed bronchial nodules | 336
mucosal hyperplasia and hypertrophy | 336
left hilar lymph nodes and tracheal nodules were biopsied | 336
TM was cultured from a bronchial nodule, left hilar lymph node, and bronchoalveolar lavage fluid | 336
NGS was performed | 336
diagnosed with disseminated TM and B. cepacia infection | 336
amphotericin B was added as antifungal therapy | 336
discontinued ceftazidime and levofloxacin | 672
cough improved | 672
febrile again | 1008
new mass appeared on the right side of the neck | 1008
chest CT scan revealed significant improvement in the pulmonary lesions | 1008
CT of the neck showed an abscess in the posterior pharyngeal wall | 1008
fracture of the 4th cervical vertebra | 1008
mass on the right side of the neck | 1008
ceftazidime and levofloxacin were added as antibacterial treatment | 1008
antibiotics were switched to meropenem and cotrimoxazole | 1056
acute-onset quadriplegia | 1104
emergency subtotal resection of the 4th cervical vertebra | 1104
widening and decompression of the spinal canal | 1104
transferred to the intensive care unit | 1104
treated with meropenem and tigecycline as antibiotics | 1104
voriconazole as an antifungal agent | 1104
B. cepacia was cultured repeatedly from the blood and pus | 1104
pulmonary lesions were improved | 1104
neck abscess could not be contained | 1104
disseminated widely to multiple body parts | 1104
hepatorenal dysfunction | 1176
cardiac insufficiency | 1176
hypotension | 1176
hypoxic | 1176
repeated immune function test | 1176
CD3+, CD4+, and CD8+ T-lymphocyte counts | 1176
disseminated intravascular coagulation | 1248
died of B. cepacia sepsis | 1248
measured the nAIGAs in the peripheral blood | 168
serum AIGA was determined by an enzyme-linked immunosorbent assay kit | 168
persistently high positive titer | 168
antibody titer increased gradually | 1344
positive titer value was based on previous study | 1344