61 years old | 0
female | 0
Caucasian | 0
admitted to the hospital | 0
peripheral arterial disease | -672
hyperlipidemia | -672
previous tobacco use | -672
midsternal chest pain | -48
acute occlusion of the right anterior artery | -2400
right common iliac artery stenting | -2400
right tibial artery stenting | -2400
stent occlusion in the right tibial artery | -672
unvaccinated for COVID-19 | 0
no respiratory symptoms | 0
no nausea | 0
no vomiting | 0
admitted to rule out acute coronary syndrome | 0
cardiology service evaluation | 0
troponins test | 0
D-dimer test | 0
vitals within normal limits | 0
heart rate in the 60s | 0
COVID-19 antigen test | 0
COVID-19 PCR test | 0
COVID-19 positive | 0
dexamethasone 6 mg IV daily | 0
NMV/r initiation | 0
apixaban 5 mg oral daily | -672
atorvastatin 40 mg oral at bedtime | -672
clopidogrel 75 mg oral daily | -672
atorvastatin held | 0
apixaban dose-adjusted to 2.5 mg twice daily | 0
nirmatrelvir 300 mg and ritonavir 100 mg twice daily | 0
heart rate decline | 12
sinus bradycardia | 24
NMV/r discontinued | 24
atropine 0.5 mg IV twice | 24
transcutaneous pacer | 24
transferred to medical ICU | 24
dobutamine drip | 24
dobutamine titrated up to 5 µg/kg/min | 24
dobutamine discontinued | 34
terbutaline tablet 5 mg by mouth | 24
terbutaline discontinued | 48
low cortisol levels | 48
cosyntropin stimulation tests | 48
MRI of the brain | 48
MRI results negative | 72
asymptomatic from COVID-19 | 120
discharged | 120