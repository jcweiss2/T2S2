85 years old | 0
female | 0
cardiac arrest | 0
cardiopulmonary resuscitation | 0
returning to spontaneous circulation | 0
urinary tract infection | -720
left pleuritic pain | -72
cough | -72
dementia | -8760
arterial hypertension | -8760
diabetes mellitus type II | -8760
depression | -8760
sedation | 0
no brain reflexes | 0
mydriatic pupils | 0
leukocytosis with neutrophilia | 0
type II myocardial infarction | 0
right basal consolidation | 0
septic shock of pulmonary origin | 0
myocardial infarction | 0
antibiotics | 0
piperacillin | 0
clarithromycin | 0
vasopressor | 0
norepinephrine | 0
mechanical ventilator support | 0
brain CT scan | 0
diffuse brain edema | 0
subfalcine herniation | 0
transtentorial herniation | 0
Glasgow Coma Scale score of 3/15 | 48
absence of brainstem reflexes | 48
brain MRI scan | 72
BOLD signal | 72
DTI acquisitions | 72
second cardiac arrest | 72
unsuccessful cardiopulmonary resuscitation | 72
death | 72
disruption of ventral and dorsal tegmental tracts | 72
reduction in FA values | 72
hyperconnective association among ARAS and cortical nuclei | 72
increased level of integration among ARAS and cortical nuclei | 72
reduction of segregation level in functions linked with consciousness | 72
breakdown of brain functional modularity | 72
abnormal propagation of information across the brain | 72
reduction of functional specialization | 72
abnormal cerebral activity | 72
admission to the hospital | 0
admission to the intensive care unit | 0
sedation withdrawal | 48
DTT demonstration of disruption of both ventral and dorsal tegmental tracts | 72
FA values computation | 72
FC estimation | 72
rsfMRI analysis | 72
DTI analysis | 72
DTT analysis | 72
neuroimaging data acquisition | -72
neuroimaging data preprocessing | 0
location and characterization of the regions of interest | 0
functional connectivity inside ARAS | 72
structural connectivity inside ARAS | 72
authorization request to Institutional Ethics Board | -72
informed consent | -72
case report review | -72
approval by Fundación Universitaria de Ciencias de la Salud Review Board | -72