79 years old | 0
female | 0
Caucasian | 0
admitted to the hospital | 0
medial femoral neck fracture | -144
low energy trauma | -144
fell on her right body side | -144
arterial hypertension | 0
hypothyreosis | 0
cataract | 0
macular degeneration | 0
hypacusis | 0
multiple operations of eyes and hand | 0
pain in her right hip | 0
abdomen presented soft | 0
no tenderness on palpation | 0
regular peristaltic sounds | 0
implanted a cemented dual head prosthesis | 24
progressive hemodynamic instability | 120
decreasing hemoglobin levels | 120
progressive serum lactate levels | 120
vasopressor-dependent | 120
intubated | 120
blood transfusion initiated | 120
free intraabdominal fluid | 120
large partially coagulated intraperitoneal hematoma | 120
free abdominal fluid | 120
suprasplenic coagulum | 120
pleural and pericardial effusion | 120
emergency splenectomy | 120
postoperative period without complications | 120
respiratory failure | 168
pneumonia | 168
septic shock | 168
multiple organ failure | 168
therapy ended | 432
died | 432
delayed splenic rupture | 120
hemorrhagic shock | 120
retroperitoneal hematoma | 120
hematoma of the thigh | 120
pseudo-aneurysms | 120
intraoperative injury | 24
branches from the common femoral artery and vein | 24
FAST-sonography not performed | 0
abdominal sonography | 120
emergency computed tomography | 120
splenectomy | 120
histopathological examination | 120
regular organ structure | 120
no preexisting splenic pathology | 0
Kehr's-sign not documented | 120
Moore stage IV | 120
large retropancreatical hematoma | 120
arterial bleeding of the pancreas | 120