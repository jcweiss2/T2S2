44 years old | 0
male | 0
Korean | 0
admitted to the hospital | 0
fever | -240
non-productive cough | -240
myalgias | -240
hypertension | -12000
treated with angiotensin-converting enzyme inhibitor | -12000
treated with oral quinolone | -168
resting dyspnea | -48
productive cough | -48
ex-smoker | 0
30-pack-a-year | 0
no history of previous respiratory diseases | 0
no specific family history | 0
temperature of 38.6℃ | 0
blood pressure of 120/80 mmHg | 0
heart rate of 90 b.p.m | 0
respiratory rate of 30 breaths/min | 0
bilateral inspiratory coarse | 0
crackles | 0
end-expiratory wheezing | 0
perihilar areas | 0
arterial blood gas values on room air | 0
pH 7.343 | 0
PaCO2 41.2 mmHg | 0
PaO2 59.2 mmHg | 0
SaO2 90.7% | 0
WBC 19,580/mm3 | 0
neutrophils 82.5% | 0
ESR 71 mm/h | 0
C-reactive protein 184.6 mg/L | 0
hemoglobin A1c 5.8% | 0
blood urea nitrogen 32.4 mg/dL | 0
creatinine 1.32 mg/dL | 0
random glucose of capillary blood 117 mg/dL | 0
bilateral bronchial wall thickening | 0
perihilar area | 0
lower lobe predominance | 0
chest X-ray | 0
sputum stains negative | 0
sputum cultures negative | 0
blood cultures negative | 0
HIV test negative | 0
empirical therapy with cefoperazone/sulbactam | 0
vancomycin | 0
high fever | 96
increasing dyspnea | 96
hypoxemia | 96
respiratory failure | 96
severe CO2 retention | 96
mechanically ventilated | 96
intensive care unit | 96
chest CT | 120
fiberoptic bronchoscopy | 120
bilateral peribronchial infiltrates | 120
patent bronchi | 120
no consolidation of the parenchyma | 120
extensive whitish exudative membranes | 120
trachea | 120
mainstem bronchi | 120
endobronchial biopsy | 120
bronchial washing fluid | 120
Aspergillus species | 120
refractory septic shock | 192
oliguria | 192
fatal cardiac arrest | 192
IV amphotericin B | 192
supportive care | 192
pseudomembranous necrotizing tracheobronchial aspergillosis | 0
invasive pulmonary aspergillosis | 0
immunocompetent host | 0
Aspergillus tracheobronchitis | 0
acute pseudomembranous tracheobronchitis | 0
Aspergillus infection | 0
tracheobronchial tree | 0
terminal respiratory failure | 192
dyspnea | -240
severe hypoxemia | 96
broad spectrum antibiotics | 0