23 years old | 0
postpartum woman | 0
septic shock | 0
transferred to the intensive care unit | 0
severe iron deficiency anemia | -672
hemoglobin concentration 8.6 g/dl | -672
gestational hypertension | -672
meconium-stained amniotic fluid | -672
prolonged rupture of the membranes | -672
chorioamnionitis | -672
urgent cesarean section | -672
developed purulent postpartum endometritis | -24
fever 39°C | -24
chills | -24
purulent uterine discharge | -24
fundal tenderness | -24
arterial line placement | -24
blood culture sample obtained | -24
initiation of empiric antibacterial therapy | -24
vancomycin | -24
gentamicin | -24
sepsis developed | -24
septic shock | -24
arterial pressure decreased to 60/40 mmHg | -24
organ failure | -24
SOFA score 16–20 | -24
Glasgow Coma Scale 10–12 points | -24
ARDS | -24
PaO2/FiO2 180 mmHg | -24
norepinephrine > 0.3 μg/kg/min | -24
bilirubin 23 mmol/L | -24
platelets 35 × 10^3/μl | -24
urine output 300 ml/day | -24
hemoglobin concentration 7.7 g/dl | -24
white blood cells 25×10^9/L | -24
prothrombin time 21 s | -24
fibrinogen concentration 89 mg/dl | -24
antithrombin III 53% | -24
D-Dimer 2.4 µg/ml | -24
C-reactive protein 309.5 mg/L | -24
procalcitonin 45 ng/ml | -24
lactate 7.5 mmol/L | -24
BNP 4,000 ng/ml | -24
normal saline bolus 30 ml/kg | -24
norepinephrine infusion 0.3 μg/kg/min | -24
intubation | -24
respiratory support assist-control mode | -24
norepinephrine increased to 3.0 μg/kg/min | -24
mean arterial pressure 60–65 mmHg | -24
mottled fingers and toes | -24
mottled abdominal wall | -24
echocardiogram showed ejection fraction 32% | -24
dobutamine infusion 20 μg/kg/min | -24
unsuccessful catecholamine dose reduction | -24
hysterectomy performed | -24
transferred to University Medical Center | -48
physical examination on admission | 0
massive aseptic necrosis of fingers I–V | 0
massive aseptic necrosis of toes I–V | 0
massive aseptic necrosis of metatarsal region | 0
massive aseptic necrosis of anterior abdominal wall | 0
sepsis/septic shock-induced multiple system failure | 0
ARDS | 0
encephalopathy | 0
systolic heart failure | 0
acute kidney injury | 0
invasive blood pressure 100/70 mmHg | 0
heart rate 150/min | 0
arterial oxygen saturation 85–92% | 0
body temperature 38.4°C | 0
sedation with dexmedetomidine | 0
mechanical ventilation assist/control | 0
PEEP 14 cmH2O | 0
FiO2 0.7 | 0
crackles over right middle and lower lung zones | 0
norepinephrine 2 μg/kg/min | 0
dobutamine 20 μg/kg/min | 0
Hb 9 g/dl | 0
WBC 22 × 10^9/L | 0
C-reactive protein 200.5 mg/L | 0
lactate 4 mmol/L | 0
procalcitonin 32 ng/ml | 0
creatine-kinase MB 15.1 IU/L | 0
BNP 5,000 ng/ml | 0
platelets 90 × 10^9/L | 0
fibrinogen 114 mg/dl | 0
activated partial thromboplastin time 128 s | 0
INR 1.27 | 0
prothrombin time 16.9 s | 0
transthoracic echocardiogram ejection fraction 38% | 0
chest radiography bilateral infiltrations | 0
PaO2/FiO2 250 mmHg | 0
blood culture Escherichia coli | 0
blood culture Pseudomonas aeruginosa | 0
blood culture Acinetobacter baumannii | 0
meropenem sensitivity | 0
no pathogens in necrotic tissues | 0
antibacterial therapy | 0
goal-directed fluid therapy | 0
nutritional support | 0
protective mechanical ventilation | 0
hydrocortisone | 0
fresh frozen plasma | 0
ascorbic acid | 0
thiamine | 0
skin wound management | 0
weaned off mechanical ventilation | 504
weaned off vasopressor therapy | 504
no neurological consequences | 504
end-organ functions returned to normal | 504
necrotic area large | 504
vasopressor support duration 8 days | 504
necrotic masses debrided | 504
autodermoplasty performed | 504
informed consent obtained | 504
23 years old|0
postpartum woman|0
septic shock|0
transferred to the intensive care unit|0
severe iron deficiency anemia|-672
hemoglobin concentration 8.6 g/dl|-672
gestational hypertension|-672
meconium-stained amniotic fluid|-672
prolonged rupture of the membranes|-672
chorioamnionitis|-672
urgent cesarean section|-672
developed purulent postpartum endometritis|-24
fever 39°C|-24
chills|-24
purulent uterine discharge|-24
fundal tenderness|-24
arterial line placement|-24
blood culture sample obtained|-24
initiation of empiric antibacterial therapy|-24
vancomycin|-24
gentamicin|-24
sepsis developed|-24
septic shock|-24
arterial pressure decreased to 60/40 mmHg|-24
organ failure|-24
SOFA score 16–20|-24
Glasgow Coma Scale 10–12 points|-24
ARDS|-24
PaO2/FiO2 180 mmHg|-24
norepinephrine > 0.3 μg/kg/min|-24
bilirubin 23 mmol/L|-24
platelets 35 × 10^3/μl|-24
urine output 300 ml/day|-24
hemoglobin concentration 7.7 g/dl|-24
white blood cells 25×10^9/L|-24
prothrombin time 21 s|-24
fibrinogen concentration 89 mg/dl|-24
antithrombin III 53%|-24
D-Dimer 2.4 µg/ml|-24
C-reactive protein 309.5 mg/L|-24
procalcitonin 45 ng/ml|-24
lactate 7.5 mmol/L|-24
BNP 4,000 ng/ml|-24
normal saline bolus 30 ml/kg|-24
norepinephrine infusion 0.3 μg/kg/min|-24
intubation|-24
respiratory support assist-control mode|-24
norepinephrine increased to 3.0 μg/kg/min|-24
mean arterial pressure 60–65 mmHg|-24
mottled fingers and toes|-24
mottled abdominal wall|-24
echocardiogram showed ejection fraction 32%|-24
dobutamine infusion 20 μg/kg/min|-24
unsuccessful catecholamine dose reduction|-24
hysterectomy performed|-24
transferred to University Medical Center|-48
physical examination on admission|0
massive aseptic necrosis of fingers I–V|0
massive aseptic necrosis of toes I–V|0
massive aseptic necrosis of metatarsal region|0
massive aseptic necrosis of anterior abdominal wall|0
sepsis/septic shock-induced multiple system failure|0
ARDS|0
encephalopathy|0
systolic heart failure|0
acute kidney injury|0
invasive blood pressure 100/70 mmHg|0
heart rate 150/min|0
arterial oxygen saturation 85–92%|0
body temperature 38.4°C|0
sedation with dexmedetomidine|0
mechanical ventilation assist/control|0
PEEP 14 cmH2O|0
FiO2 0.7|0
crackles over right middle and lower lung zones|0
norepinephrine 2 μg/kg/min|0
dobutamine 20 μg/kg/min|0
Hb 9 g/dl|0
WBC 22 × 10^9/L|0
C-reactive protein 200.5 mg/L|0
lactate 4 mmol/L|0
procalcitonin 32 ng/ml|0
creatine-kinase MB 15.1 IU/L|0
BNP 5,000 ng/ml|0
platelets 90 × 10^9/L|0
fibrinogen 114 mg/dl|0
activated partial thromboplastin time 128 s|0
INR 1.27|0
prothrombin time 16.9 s|0
transthoracic echocardiogram ejection fraction 38%|0
chest radiography bilateral infiltrations|0
PaO2/FiO2 250 mmHg|0
blood culture Escherichia coli|0
blood culture Pseudomonas aeruginosa|0
blood culture Acinetobacter baumannii|0
meropenem sensitivity|0
no pathogens in necrotic tissues|0
antibacterial therapy|0
goal-directed fluid therapy|0
nutritional support|0
protective mechanical ventilation|0
hydrocortisone|0
fresh frozen plasma|0
ascorbic acid|0
thiamine|0
skin wound management|0
weaned off mechanical ventilation|504
weaned off vasopressor therapy|504
no neurological consequences|504
end-organ functions returned to normal|504
necrotic area large|504
vasopressor support duration 8 days|504
necrotic masses debrided|504
autodermoplasty performed|504
informed consent obtained|504
