58 years old | 0
woman | 0
presented to the emergency department | 0
progressive lumbar back pain | -504
radiating to left leg | -504
sensation of numbness in lower left leg and foot | -504
symptoms progressing for past 3 weeks | -504
gait disorder | -120
lack of coordination in left foot | -120
urine incontinence | -120
bowel incontinence | -120
no abdominal pain | 0
fever 1 day prior to complaints | -24
weight loss of 11 kg | -720
appeared ill | 0
body temperature of 38.8°C | 0
decreased strength in left leg | 0
positive Lasègue sign on left side | 0
soft abdomen | 0
non-tender abdomen | 0
leukocytosis | 0
elevated C-reactive protein | 0
urine retention of 1,300 ml | 0
worsened septic condition | 0
high-grade fever (40.9°C) | 0
started Amoxicillin/Clavulanate | 0
transferred to intensive care unit | 0
MRI showing fistula from sigmoid colon to presacral abscess | 0
abscess expanded into spinal canal | 0
sacral osteomyelitis | 0
diffuse meningeal staining of conus medullaris and cauda equina | 0
chest/abdominal CT scan showing pleural fluid | 0
multiple fluid and air collections | 0
air in spinal canal and back muscles | 0
Hartmann's procedure performed | 0
intra-abdominal abscesses drained | 0
intra-abdominal drains placed | 0
postoperative management with broad-spectrum antibiotics | 0
therapeutic heparin for thrombus in left iliac vein | 0
extubated on postoperative day one | 24
transferred to gastrointestinal surgery ward on postoperative day four | 96
stoma production started | 96
persisting neurological symptoms | 336
returned to primary care center | 336
enrolled in intensive rehabilitation program | 336
cauda equina syndrome | 0
fistula formation to spinal cord | 0
complicated diverticulitis | 0
pelvic abscess | 0
purulent peritonitis | 0
thrombus in left iliac vein | 0
hemodynamically normal | 0
no signs of spondylodiscitis | 0
no abnormalities on chest and lumbar spine X-ray | 0
unable to urinate initially | 0
denied abdominal pain | 0
denied chest pain | 0
denies shortness of breath | 0
no rectal device mentioned | 0
normal sensation in saddle area | 0
normal perianal area | 0
normal anal sphincter tone | 0
no epidural abscess | 0
no colon cancer | 0
no spondylodiscitis | 0
no fecal peritonitis | 0
no intestinal obstruction | 0
no colovesical fistula | 0
no colovaginal fistula | 0
no coloenteric fistula | 0
no colocutaneous fistula | 0
no involvement of intervertebral discs | 0
no emergency surgery indicated initially | 0
no primary anastomosis made | 0
no complete resolution of neurological symptoms | 0
no significant pain postoperatively | 0
no signs of sepsis postoperatively | 0
no recurrence of abscess | 0
no postoperative infection | 0
no complications during rehabilitation | 0
no further weight loss postoperatively | 0
no evidence of colon cancer | 0
no urinary tract infection | 0
no respiratory complications | 0
no hemodynamic instability postoperatively | 0
no signs of wound infection | 0
no evidence of recurrent diverticulitis | 0
no further episodes of incontinence postoperatively | 0
no recurrence of fever postoperatively | 0
no further episodes of urinary retention | 0
no signs of heparin-induced thrombocytopenia | 0
no allergic reactions to antibiotics | 0
no adverse drug reactions | 0
no postoperative bleeding | 0
no anastomotic leak | 0
no stoma complications | 0
no evidence of venous thromboembolism post-thrombus | 0
no recurrence of thrombus | 0
no further episodes of cauda equina syndrome | 0
no complications during intensive rehabilitation | 0
no further episodes of back pain | 0
no recurrence of numbness | 0
no further gait disorder | 0
no signs of recurrent osteomyelitis | 0
no further meningeal staining | 0
no recurrence of presacral abscess | 0
no further fluid collections postoperatively | 0
no recurrence of air in spinal canal | 0
no evidence of recurrent fistula | 0
no postoperative ileus | 0
no evidence of malnutrition | 0
no evidence of dehydration | 0
no electrolyte imbalances postoperatively | 0
no evidence of anemia postoperatively | 0
no evidence of thrombocytopenia | 0
no evidence of leukopenia | 0
no signs of adrenal insufficiency | 0
no evidence of hypothyroidism | 0
no evidence of liver dysfunction | 0
no evidence of renal dysfunction postoperatively | 0
no evidence of pancreatitis | 0
no evidence of diabetes mellitus | 0
no evidence of glucose intolerance | 0
no evidence of coagulopathy beyond INR elevation | 0
no evidence of hyperglycemia requiring insulin | 0
no evidence of hypokalemia | 0
no evidence of hyponatremia | 0
no evidence of hypercalcemia | 0
no evidence of hypomagnesemia | 0
no evidence of hypophosphatemia | 0
no evidence of hypozincemia | 0
no evidence of vitamin deficiencies | 0
no evidence of trace element deficiencies | 0
no evidence of protein-energy malnutrition | 0
no evidence of overhydration | 0
no evidence of fluid overload | 0
no evidence of heart failure | 0
no evidence of arrhythmias | 0
no evidence of myocardial infarction | 0
no evidence of pericarditis | 0
no evidence of endocarditis | 0
no evidence of pulmonary embolism | 0
no evidence of pneumonia | 0
no evidence of asthma exacerbation | 0
no evidence of COPD exacerbation | 0
no evidence of allergic rhinitis | 0
no evidence of sinusitis | 0
no evidence of otitis media | 0
no evidence of pharyngitis | 0
no evidence of tonsillitis | 0
no evidence of gastroenteritis | 0
no evidence of food poisoning | 0
no evidence of hepatitis | 0
no evidence of cholecystitis | 0
no evidence of appendicitis | 0
no evidence of peptic ulcer disease | 0
no evidence of gastritis | 0
no evidence of esophagitis | 0
no evidence of inflammatory bowel disease | 0
no evidence of celiac disease | 0
no evidence of lactose intolerance | 0
no evidence of food allergies | 0
no evidence of autoimmune disorders | 0
no evidence of rheumatoid arthritis | 0
no evidence of lupus | 0
no evidence of vasculitis | 0
no evidence of sarcoidosis | 0
no evidence of amyloidosis | 0
no evidence of hemochromatosis | 0
no evidence of porphyria | 0
no evidence of connective tissue disorders | 0
no evidence of Marfan syndrome | 0
no evidence of Ehlers-Danlos syndrome | 0
no evidence of neurofibromatosis | 0
no evidence of tuberous sclerosis | 0
no evidence of Huntington's disease | 0
no evidence of Parkinson's disease | 0
no evidence of multiple sclerosis | 0
no evidence of Guillain-Barré syndrome | 0
no evidence of myasthenia gravis | 0
no evidence of ALS | 0
no evidence of dementia | 0
no evidence of delirium | 0
no evidence of psychosis | 0
no evidence of depression | 0
no evidence of anxiety | 0
no evidence of bipolar disorder | 0
no evidence of schizophrenia | 0
no evidence of personality disorders | 0
no evidence of eating disorders | 0
no evidence of substance abuse | 0
no evidence of alcohol use disorder | 0
no evidence of nicotine dependence | 0
no evidence of opioid dependence | 0
no evidence of stimulant use disorder | 0
no evidence of cannabis use disorder | 0
no evidence of hallucinogen use disorder | 0
no evidence of gambling disorder | 0
no evidence of internet addiction | 0
no evidence of gaming disorder | 0
no evidence of sex addiction | 0
no evidence of other behavioral addictions | 0
no evidence of sleep disorders | 0
no evidence of insomnia | 0
no evidence of sleep apnea | 0
no evidence of narcolepsy | 0
no evidence of circadian rhythm disorders | 0
no evidence of parasomnias | 0
no evidence of movement disorders | 0
no evidence of restless leg syndrome | 0
no evidence of tic disorders | 0
no evidence of Tourette syndrome | 0
no evidence of dystonia | 0
no evidence of chorea | 0
no evidence of ataxia | 0
no evidence of vertigo | 0
no evidence of Meniere's disease | 0
no evidence of labyrinthitis | 0
no evidence of benign positional vertigo | 0
no evidence of vestibular neuritis | 0
no evidence of acoustic neuroma | 0
no evidence of hearing loss | 0
no evidence of tinnitus | 0
no evidence of visual disturbances | 0
no evidence of glaucoma | 0
no evidence of cataracts | 0
no evidence of macular degeneration | 0
no evidence of diabetic retinopathy | 0
no evidence of hypertensive retinopathy | 0
no evidence of uveitis | 0
no evidence of keratitis | 0
no evidence of conjunctivitis | 0
no evidence of blepharitis | 0
no evidence of orbital cellulitis | 0
no evidence of optic neuritis | 0
no evidence of papilledema | 0
no evidence of corneal abrasion | 0
no evidence of dry eye syndrome | 0
no evidence of allergic conjunctivitis | 0
no evidence of seasonal allergies | 0
no evidence of perennial allergies | 0
no evidence of atopic dermatitis | 0
no evidence of contact dermatitis | 0
no evidence of psoriasis | 0
no evidence of eczema | 0
no evidence of urticaria | 0
no evidence of acne | 0
no evidence of rosacea | 0
no evidence of vitiligo | 0
no evidence of alopecia | 0
no evidence of fungal infections | 0
no evidence of bacterial infections | 0
no evidence of viral infections | 0
no evidence of parasitic infections | 0
no evidence of scabies | 0
no evidence of lice infestation | 0
no evidence of cellulitis | 0
no evidence of erysipelas | 0
no evidence of impetigo | 0
no evidence of folliculitis | 0
no evidence of necrotizing fasciitis | 0
no evidence of Stevens-Johnson syndrome | 0
no evidence of toxic epidermal necrolysis | 0
no evidence of drug eruptions | 0
no evidence of erythema multiforme | 0
no evidence of pemphigus | 0
no evidence of pemphigoid | 0
no evidence of bullous dermatoses | 0
no evidence of cutaneous lymphoma | 0
no evidence of melanoma | 0
no evidence of basal cell carcinoma | 0
no evidence of squamous cell carcinoma | 0
no evidence of actinic keratosis | 0
no evidence of seborrheic keratosis | 0
no evidence of molluscum contagiosum | 0
no evidence of warts | 0
no evidence of herpes simplex | 0
no evidence of herpes zoster | 0
no evidence of Lyme disease | 0
no evidence of syphilis | 0
no evidence of tuberculosis | 0
no evidence of leprosy | 0
no evidence of histoplasmosis | 0
no evidence of coccidioidomycosis | 0
no evidence of blastomycosis | 0
no evidence of cryptococcosis | 0
no evidence of aspergillosis | 0
no evidence of mucormycosis | 0
no evidence of candidiasis | 0
no evidence of pneumocystis pneumonia | 0
no evidence of toxoplasmosis | 0
no evidence of malaria | 0
no evidence of dengue fever | 0
no evidence of yellow fever | 0
no evidence of Zika virus | 0
no evidence of Ebola virus | 0
no evidence of Marburg virus | 0
no evidence of Lassa fever | 0
no evidence of rabies | 0
no evidence of tetanus | 0
no evidence of diphtheria | 0
no evidence of pertussis | 0
no evidence of measles | 0
no evidence of mumps | 0
no evidence of rubella | 0
no evidence of chickenpox | 0
no evidence of scarlet fever | 0
no evidence of rheumatic fever | 0
no evidence of Kawasaki disease |;end of text|>
