66 years old | 0
male | 0
T1 high grade transitional cell carcinoma of a bladder diverticulum | -672
radical cystoprostatectomy | 0
ileal conduit formation | 0
lobectomy for primary lung adenocarcinoma | -10080
sigmoid colectomy for stage II colon adenocarcinoma | -10080
type 2 diabetes | 0
hypertension | 0
previous cardiac stenting | 0
high grade small bowel obstruction | 120
exploratory laparotomy | 120
interstitial herniation of small bowel | 120
aspiration of gastric contents | 120
difficulties with ventilation | 120
oxygenation | 120
sepsis | 120
venous-venous extracorporeal membrane oxygenation | 120
weaned off VV-ECMO | 240
extubated | 240
septic shock | 240
vasopressor requirements increasing | 240
inotropic requirements increasing | 240
computed tomography scan of the abdomen | 240
new widespread free fluid | 240
bowel oedema | 240
new ischaemic bowel | 240
small anastomotic leak | 240
Hartmann's resection | 240
anastomotic leak managed conservatively | 240
Bander ureteral diversion stents | 240
persistent uretero-ileal anastomotic leaks | 480
ongoing sepsis | 480
vasopressor requirements | 480
new pelvic collection | 480
urethral indwelling catheter | 480
Flexi-Seal rectal tube | 480
free drainage of the pelvic collection | 480
creatinine level | 480
urinary diversion with bilateral nephrostomy tubes | 720
persistent leak from uretero-ileal anastomosis | 720
methylene blue injection | 720
nephrostograms | 720
free drainage into the pelvic collection | 720
ureteric embolisation | 720
Interlock-18 coils | 720
Histoacryl/Lipiodol glue | 720
satisfactory occlusion | 720
covering 10.2Fr nephrostomy tube | 720
repeat nephrostogram | 1008
ongoing leak beyond the right embolisation coil | 1008
ongoing sepsis | 1008
another attempt at embolisation | 1008
MVP-9Q plug | 1008
Histoacryl/Lipiodol in 1:3 dilution | 1008
final nephrostogram | 1008
adequate occlusion of the ureters | 1008
transferred to a rehabilitation facility | 1344
bilateral nephrostomy tubes | 1344
all other drains and tubes removed | 1344
discharged home | 1344
ongoing follow-up with the Urology service | 1344
regular 6-weekly nephrostomy tube exchanges | 1344
nephrostogram to assess embolisation site | 1344
surveillance scans for bladder cancer | 1344