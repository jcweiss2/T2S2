86 years old | 0  
    male | 0  
    chronic heart failure | 0  
    atrial fibrillation | 0  
    followed by a cardiologist as an outpatient | 0  
    admitted to the ICU | 0  
    septic shock | 0  
    urinary tract infection | 0  
    Charlson morbidity score of 7 | 0  
    respiratory distress | 0  
    required intubation | 0  
    mechanical ventilation | 0  
    advanced care preferred | 0  
    impaired level of consciousness | 0  
    consent from family for life-sustaining therapy | 0  
    antibiotic therapy | 0  
    management of mechanical ventilation | 0  
    physical status recovered temporarily | 0  
    reduction in level of consciousness | -864  
    brain infarction | -864  
    informed family of poor prognosis | -864  
    acute panperitonitis | -1152  
    gastrointestinal perforation | -1152  
    proposed operation or conservative care | -1152  
    family selected conservative management | -1152  
    physical condition worsened | -1176  
    oliguria | -1176  
    progression of renal insufficiency | -1176  
    consulted nephrologists | -1176  
    hemodialysis proposed | -1176  
    systolic blood pressure maintained at 80 mm Hg | -1176  
    continuous intravenous vasopressor | -1176  
    uncontrollable sepsis | -1176  
    multiple organ failure | -1176  
    marked thrombocytopenia | -1176  
    insertion of dialysis catheter risk | -1176  
    discussed with cardiologists, nephrologists, nurses | -1176  
    concluded HD not effective or safe | -1176  
    recognized palliative care as acceptable | -1176  
    explained HD not beneficial | -1176  
    referred to palliative care (NTD) | -1176  
    family withheld decision | -1176  
    family agreed to NTD | -1200  
    patient died | -1248  
    family satisfied with care | -1248  

