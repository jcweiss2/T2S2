75 years old | 0
female | 0
visited emergency room | 0
dyspnea | -168
idiopathic thrombocytopenic purpura | -720
corticosteroids | -720
prednisolone | -720
admitted to intensive care unit | 0
empirical treatment | 0
community-acquired pneumonia | 0
intravenous piperacillin/tazobactam | 0
azithromycin | 0
IV sulfamethoxazole/trimethoprim | 0
methylprednisolone | 0
endotracheal intubation | 72
mechanical ventilator support | 72
antibiotics switched to meropenem | 72
levofloxacin | 72
fraction of inspiration O2 reduced | 168
clinical improvement | 168
initial serology | 168
PCP PCR positive | 168
aspergillus antigen positive | 168
itraconazole | 168
follow-up non-enhanced chest CT | 168
newly formed GGOs | 168
cavitary changes | 168
bedside bronchoscopy | 216
bronchoalveolar lavage | 216
PCP PCR | 216
aspergillus antigen | 216
aspergillosis reported | 264
IA diagnosed | 264
antifungal agent changed to voriconazole | 264
percutaneous dilatational tracheostomy | 312
bronchoscopy with BAL | 312
BAL fluid cytology | 312
condition deteriorated | 360
family declined aggressive management | 360
extracorporeal membrane oxygenation declined | 360
PCP PCR of BAL fluid specimen positive | 360
fungus culture no growth | 360
multi-organ failure | 384
septic shock | 384
died | 384