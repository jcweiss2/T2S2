23 years old | 0
male | 0
admitted to the hospital | 0
abdominal pain | 0
nausea | 0
vomiting | 0
diarrhea | 0
pulseless electrical activity cardiac arrest | 0
peripheral venoarterial ECMO | 0
healthy individual | -672
no past medical history | -672
septic shock | 0
hypovolemic shock | 0
cardiovascular failure | 0
transthoracic echocardiogram | 0
near cardiac standstill | 0
moderate posterior pericardial effusion | 0
systolic blood pressure 30 mm Hg | 0
low ECMO flow | 0
bridge circuit | 0
no change in flow | 0
augment venous drainage | 0
right internal jugular venous cannula | 0
venovenous-arterial ECMO | 0
blood pressure improved | 0
increased venous drainage | 0
better ECMO flow | 0
hemodynamically unstable | 0
pericardial effusion enlarged | 0
emergent pericardiotomy | 0
400 ml clear fluid removed | 0
severe myocardial edema | 0
near cardiac standstill | 0
left ventricle nonpulsatile | 0
competing with retrograde ECMO flow | 0
severe LV dilation | 0
pulmonary edema | 0
Impella CP heart pump placement | 0
LV venting | 0
opening aortic pressure 72/64 mm Hg | 0
LV end-diastolic pressure 25 mm Hg | 0
LV cavity size decreased | 0
improved unloading from Impella CP | 0
lower extremities became tense | 0
creatinine kinase level rose | 0
severe fulminant skeletal myositis | 0
H3N2 viremia | 0
rhabdomyolysis | 0
bilateral leg fasciotomies | 0
removal of Impella device | 0
oseltamivir treatment | 0
broad-spectrum antibiotics | 0
respiratory swab positive for influenza A | 0
blood cultures grew Streptococcus viridans | 0
fulminant myocarditis | 0
intravenous immunoglobulin | 0
ECMO flow requirement decreased | 24
cardiac contractility increased | 24
TTE on hospital day 12 | 288
estimated LV ejection fraction 30-35% | 288
lungs severely damaged | 288
differential upper extremity hypoxemia | 288
North-South syndrome | 288
ECMO circuit rearranged | 288
VA-venous configuration | 288
oxygenated blood returned to upper body | 288
improved oxygenation | 288
facial swelling | 288
superior vena cava syndrome | 288
cannula removed | 288
facial swelling resolved | 288
ECMO configuration switched | 288
VA through left femoral artery and vein | 288
hemodynamic improvement | 288
vasopressor requirements decreased | 432
ECMO circuit decannulated | 432
multiple infections | 432
extensive wound debridement | 432
tracheostomy placed | 432
tracheostomy decannulated | 432
weaned off hemodialysis | 432
TTE showed LV ejection fraction 55% | 432
discharged | 432