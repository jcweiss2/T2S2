50 years old | 0
male | 0
admitted to the hospital | 0
chronic pancreatitis | 0
chronic alcohol use | -17280
epigastric abdominal pain | -1440
generalized weakness | -1440
chronic abdominal pain | -17280
denied nausea | 0
denied vomiting | 0
denied diarrhea | 0
denied constipation | 0
denied change in urinary habits | 0
denied recent travel | 0
denied sick contacts | 0
acetaminophen | -17280
oxycodone | -17280
pancreatic enzyme replacement therapy | -17280
blood pressure 100/92 mm Hg | 0
heart rate 94 bpm | 0
respiratory rate 16 breaths/min | 0
O2 saturation 97% | 0
epigastric tenderness | 0
computed tomography abdomen | -17280
pancreas with diffuse calcifications | -17280
hyperglycemic | 0
blood glucose 703 mg/dL | 0
serum bicarbonate 16 mmol/L | 0
ketones in urine | 0
acetone in blood | 0
anion gap corrected for albumin 27 | 0
DKA | 0
admitted to medical intensive care unit | 0
nil per os | 0
intravenous lactated Ringer's solution | 0
potassium | 0
IV insulin drip | 0
pancreatic enzyme replacement held | 0
cardiac enzymes sent | 0
lipase sent | 0
cardiac enzymes normal | 0
lipase elevated 156 | 0
septic workup sent | 0
septic workup negative | 0
blood glucose monitored every hour | 0
electrolytes monitored every 4 hours | 0
albumin monitored every 4 hours | 0
IV hydration continued | 0
adjustments of potassium | 0
adjustments of dextrose | 0
anion gap closed | 0
transitioned to insulin detemir 10 Units SQ QHS | 0
diabetic diet 2 hours after detemir | 0
insulin sliding scale | 0
sent to medical floor | 0
diabetic teaching provided | 0
insulin regimen optimized | 0
discharged | 0
insulin aspart 3 Units TID | 0
insulin detemir 10 Units QHS | 0
insulin detemir 6 Units QAM | 0
autoimmune workup sent | 0
autoimmune workup negative | 0
ketorolac for abdominal pain | 0
follow up with primary care physician | 0
prior HbA1c normal | -17280
HbA1c 16% | 0
DM3c diagnosis | 0
DKA presentation | 0
