34 years old | 0
male | 0
Marfan syndrome | 0
Bentall procedure in 2018 | -17520
admitted with worsening dyspnea (NYHA class IV) | 0
tachycardia | 0
fever | 0
suspected infective endocarditis | 0
heart rate 118 beats/min | 0
blood pressure 92/45 mmHg | 0
peripheral oxygen saturation 85% | 0
body temperature 38.6°C | 0
COVID-19 positive | 0
moved to negative-pressure ICU room | 0
bilateral ground glass opacities | 0
interlobular septal thickening | 0
dependent consolidation | 0
mechanical bileaflet prosthetic valve | 0
suspected vegetations on the leaflets | 0
dehiscence of the aortic root | 0
para-aortic abscess | 0
moderate aortic regurgitation | 0
no pericardial effusion | 0
contrast leakage in mediastinum | 0
normal ascending aorta, arch, and descending aorta | 0
anemia | 0
leukocytosis |! 0
thrombocytopenia | 0
high procalcitonin | 0
high interleukin-6 | 0
bacterial cultures negative | 0
meropenem started | 0
vancomycin started | 0
remdesivir infusion (loading dose 200 mg IV) | 0
remdesivir (100 mg once/day) | 0
urgent cardiac surgery advised | 0
EuroSCORE II 10.82% | 0
redo Bentall surgery in negative-pressure operating room | 0
invasive arterial pressure monitoring | 0
pulmonary artery catheter | 0
transesophageal echocardiography | 0
cerebral oximetry | 0
cardiopulmonary bypass instituted | 0
axillary artery cannulation | 0
femoral vein cannulation | 0
moderate hypothermia | 0
Custodiol cardioplegia | 0
alpha-stat blood gas management | 0
CytoSorb hemoadsorber integrated into CPB circuit | 0
CytoSorb used for entire CPB duration | 0
redo sternotomy | 0
cleaning para-aortic pus | 0
extraction of previous valve graft | 0
creation of neo-annulus with bovine pericardium | 0
redo Bentall procedure with porcine root | 0
no infective endocarditis intraoperatively | 0
aortic-cross clamp time 165 min | 0
cardiopulmonary bypass duration 191 min | 0
epinephrine 0.05 µg/kg/min | 0
norepinephrine 0.3 µg/kg/min | 0
red blood cells transfusion (10 units) | 0
fresh frozen plasma transfusion (6 units) | 0
platelet apheresis transfusion (4 units) | 0
excessive bleeding | 0
pre-existing anemia | 0
pre-existing thrombocytopenia | 0
transferred back to ICU | 0
weaned from ventilator after 48 hours | 48
weaned from inotropes after 48 hours | 48
inflammatory markers improved postoperatively | 48
hemodynamic parameters improved postoperatively | 48
uneventful remaining hospital stay | 48
Bentall procedure in 2018 | -26280
leukocytosis | 0
