1-year-old| 0
male | 0
presented to Accident and Emergency department | 0
irritable | 0
drowsy | 0
Glasgow Coma Score 7 | 0
mild right-sided weakness | 0
unequal pupils | 0
right pupil 5+ | 0
left pupil 3+ | 0
no external injuries | 0
intra-osseous needle placed in right tibia | 0
intubated | 0
induction with fentanyl 2 mcg/kg | 0
induction with propofol 2 mg/kg | 0
induction with rocuronium 0.8 mg/kg | 0
hand ventilated | 0
maintained normal end-tidal carbon dioxide | 0
head computed tomography scan | 0
acute right-sided subdural hematoma | 0
significant midline shift | 0
transferred to operating theater | 0
right frontal craniotomy | 0
evacuation of acute subdural hematoma | 0
systolic blood pressure 98 mmHg | 0
good pulses | 0
mottled peripheries | 0
pale blue skin | 0
venous access through left femoral triple lumen central line | 0
arterial pressure monitoring through right femoral 22G cannula | 0
tympanic membrane temperature 36.0°C | 0
received 30 ml/kg 3% hypertonic saline | 0
surgery commenced | 0
anesthesia maintained with O2/N2O | 0
anesthesia maintained with sevoflurane | 0
positive pressure ventilation | 0
large volume of urine passed | 0
Hartmann's solution 400 ml infused | 0
Hartmann's solution in 5 ml/kg boluses | 0
maintained blood pressure during anesthesia | 0
moderate blood loss | 0
transfusion not required | 0
arterial blood gas during surgery | 0
mixed respiratory acidosis | 0
pH 7.08 | 0
PCO2 9.2 KPa | 0
PO2 31.6 KPa | 0
Na+ 154 mmol/L | 0
K+ 3.0 mmol/L | 0
Cl 129 mmol/L | 0
Ca++ 1.36 mmol/L | 0
glucose 14.1 mmol/L | 0
lactate 0.8 mmol/L | 0
hemoglobin 10.0 g/L | 0
base excess -9.8 | 0
highest serum sodium 158 mmol/L | 0
hemoglobin 8.0 g/dl at end of surgery | 0
right fronto2-occipital hematoma evacuated | 0
transported to pediatric Intensive Care Unit | 0
ventilated | 0
sedated with midazolam 3 mcg/kg/min | 0
sedated with morphine 20 mcg/kg/h | 0
extubated 2 hours after surgery | 24
postoperative fluid intake 2/3rd of daily requirement orally | 24
good urine output 1-2 ml/kg/h | 24
SaO2 98%-100% | 24
self-ventilating room air | 24
respiratory rate 24-28 bpm | 24
no respiratory distress | 24
heart rate 140/min | 24
blood pressure 112/66 mmHg | 24
pupils equal | 24
pupils reacted to light | 24
awake | 24
alert | 24
electrolytes normal Na+ 139-141 mmol/L | 24
lower and normalizing K+ 3.4-3.8 mmol/L | 24
temperature spike 38.8°C | 24
temperature spike resolved with paracetamol | 24
drug error explained to parents | 24
uneventful recovery | 24
no detectable residual defects | 24
no renal injury | 24
no residual brain damage | 24
normal electrolytes at follow-up after 1 month | 720
