59 years old | 0
female | 0
admitted to the hospital | 0
high temperature | 0
orthostatic hypotension | 0
left thigh pain | 0
back pain | -360
fever | -48
chills | -48
sweats | -48
extreme fatigue | -48
antipyretic agents | -48
temperature rose to 39.5 °C | -24
unbearable thigh pain | -24
surgical procedure to the left ilium | -47520
staphylococcal osteomyelitis | -47520
hypotension | 0
systolic pressure of 70 mmHg | 0
pulse of 90 beats per minute | 0
normal temperature | 0
respiratory rate of 15 breaths per minute | 0
oxygen saturation of 96% | 0
thigh sensitivity | 0
pain to the left hip and thigh | 0
mildly elevated white blood cell count | 0
neutrophilic predominance | 0
elevated inflammatory markers | 0
mildly elevated liver enzymes | 0
elevated creatinine kinase | 0
febrile | 0
blood cultures | 0
antipyretics | 0
empirical antibiotics | 0
abscess within the left iliopsoas muscle | 0
abscesses in the gluteus muscle | 0
CT guidance | 0
pus aspiration | 0
new-onset sudden bilateral pleuritic pain | 12
difficulty in breathing | 12
abnormal breath sounds | 12
crackles | 12
diffuse rhonchi | 12
hypoxia | 12
bilateral opacities | 12
nodular infiltrates in both pulmonary fields | 12
septic pulmonary emboli | 12
acute respiratory distress syndrome | 12
right-sided endocarditis | 12
thrombosis in the lower extremities | 12
mechanical ventilation | 24
methicillin-susceptible strain of S. aureus | 120
linezolid 600 mg intravenously | 120
weaned from the ventilator | 168
repeated CT | 360
reduction of the iliopsoas abscess | 360
cavitation of the nodular lung infiltrates | 360
intravenous antibiotics | 720
oral treatment | 1440
repeated CT | 2160
complete disappearance of abscesses | 2160