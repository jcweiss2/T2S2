30 years old | 0
male | 0
end-stage renal disease | -672
hypertensive nephropathy | -672
renal transplant | -128
deceased-donor kidney transplant | -128
tacrolimus | -128
mycophenolate mofetil | -128
prednisone acetate | -128
metoprolol succinate | -128
generalized pain | -72
headache | -72
fever | -72
palpitation | -72
watery diarrhea | -24
poor mental status | 0
highest temperature of 38.4 ℃ | 0
blood pressure reading of 80/60 mmHg | 0
leukocyte count of 10.38×10^9/L | 0
neutrophil percentage of 90% | 0
hemoglobin of 63 g/L | 0
serum creatinine level of 344 µmol/L | 0
infusions of suspended red blood cells | 0
CMV infection | -128
BK virus infection | -128
graft rejection | -128
intravenous cefoperazone sulbactam | 24
convulsions | 144
headaches | 144
diplopia | 144
meningeal irritation sign negative | 144
maximum body temperature of 40.0 ℃ | 144
pulse rate of 64–120 beats/min | 144
respiratory rate of 16–39 breaths/min | 144
white blood cell count of 5.34×10^9/L | 144
neutrophil percentage of 92% | 144
procalcitonin of 3.2 mg/L | 144
total protein of 2.37 g/L | 144
chloride of 125.3 mmol/L | 144
glucose of 4.36 mmol/L | 144
Lm detected in blood culture | 144
Lm detected in cerebrospinal fluid culture | 216
cranial MRI scan | 192
lesions in the posterior horn of the left lateral ventricle | 192
sodium penicillin infusion pump | 216
levetiracetam tablets | 216
methylprednisolone | 216
FK-506 discontinued | 216
MMF discontinued | 216
allergic reaction to penicillin | 240
rashes on lower back and four limbs | 240
compound sulfamethoxazole tablets | 240
TMP-SMX 960 mg every 6 hours | 240
tracheal intubation removed | 408
oral treatment with TMP-SMX 960 mg every 12 hours | 408
immunosuppressant therapy resumed | 408
temperature of 36.7 ℃ | 528
hemoglobin level of 83 g/L | 528
white blood cell count of 4.51×10^9/L | 528
neutrophil percentage of 72.4% | 528
CSF yellowish and protein-negative | 528
chlorine of 123.6 mmol/L | 528
glucose of 123.6 mmol/L | 528
SCr of 269.8 µmol/L | 528
T2 hyperdense shadow in the brain | 528
cranial MRI 6 months after discharge | 1056
gliosis smaller | 1056
absorption of mastoiditis smaller | 1056