75 years old | 0
    woman | 0
    presented at the accident and emergency department | 0
    epigastric pain | -48
    right upper quadrant pain | -48
    nausea | -48
    no fever | -48
    referred for nonspecific digestive difficulties | -2016
    similar episode 1 week earlier | -168
    unremarkable cardiorespiratory examination | 0
    hemodynamically stable | 0
    tender abdomen | 0
    guarding in the right upper quadrant | 0
    positive Murphy's sign | 0
    gallbladder distension | 0
    gallbladder wall thickening | 0
    2.5 cm stone in the gallbladder lumen | 0
    no pericholecystic fluid | 0
    no intrahepatic ductal dilatation | 0
    no extrahepatic ductal dilatation | 0
    white blood cell count 8.3 × 10^9/l | 0
    C-reactive protein 85 mg/l | 0
    serum total bilirubin 17.3 µmol/l | 0
    alkaline phosphatase 79 IU/l | 0
    aspartate aminotransferase 23 IU/l | 0
    alanine aminotransferase 29 IU/l | 0
    lipase 32 IU/l | 0
    sodium 136 mmol/l | 0
    potassium 3.8 mmol/l | 0
    blood urea 5.1 mmol/l | 0
    creatinine 82 µmol/l | 0
    troponin I <0.01 U/l | 0
    acute cholecystitis diagnosis | 0
    sinus rhythm | 0
    incomplete right branch block | 0
    negative T waves in V1–V3 | 0
    no sign of ischemia | 0
    intravenous antibiotics | 0
    cephalosporin | 0
    metronidazole | 0
    fluids administration | 0
    fever (39°C) | 24
    two peripheral blood cultures taken | 24
    negative blood cultures | 24
    increased white blood cell count (10.2 × 10^9/l) | 24
    CRP 434 mg/l | 24
    normal urea | 24
    normal electrolytes | 24
    normal liver function | 24
    normal amylase | 24
    normal bilirubin | 24
    surgical cholecystectomy planned | 24
    no chest pain | 24
    further preoperative ECG performed | 24
    ST segment depression in V3 | 24
    negative T waves in V1–V3 | 24
    troponin I level elevated (0.78 μg/l) | 24
    creatine kinase level 409 U/l | 24
    anticoagulation with high-dose low-molecular-weight heparin | 24
    aspirin | 24
    β-blockers | 24
    angiotensin-converting enzyme inhibitors | 24
    admitted to the intensive care unit | 24
    troponin level decreased to 0.49 μg/l after 12 hours | 36
    troponin level decreased to 0.30 μg/l after another 8 hours | 44
    mildly enlarged right ventricle | 24
    no enlargement of the left ventricle | 24
    good ejection fraction | 24
    right overload septal motion abnormality | 24
    pulmonary hypertension (systolic peripheral arterial pressure ∼45–50 mm Hg) | 24
    angio-CT performed to exclude pulmonary embolism | 24
    negative angio-CT findings | 24
    coronary angiography undertaken | 24
    no abnormality | 24
    normal left ventricular function | 24
    abdominal CT confirmed cholecystitis | 24
    excluded empyema | 24
    excluded abscess complications | 24
    progressive disappearance of abdominal symptoms | 24
    return to normal complete blood count | 24
    return to normal lipase | 24
    return to normal cardiac markers | 24
    return to normal electrolytes | 24
    return to normal bilirubin | 24
    return to normal aminotransferase | 24
    return to normal CRP levels | 24
    discharged | 24
    elective surgery for symptomatic cholelithiasis planned | 24
    <|eot_id|>
    