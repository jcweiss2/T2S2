61 years old | 0
female | 0
general weakness | -72
fall at home | -72
infected heel pressure ulcer | -72
admitted to the Department of General Surgery | 0
urinary tract infection | 0
thyroid dysfunction | 0
hemodynamic instability | 6
loss of consciousness | 6
admitted to the ICU | 6
intubated | 6
unconscious | 6
hypothermic | 6
hemodynamically unstable | 6
hypotensive | 6
bradycardic | 6
obese | 6
generalized subcutaneous edema | 6
macerated skin | 6
extensive heel pressure ulcer | 6
soft abdomen | 6
inaudible peristalsis | 6
irreducible ventral hernia | 6
hypercapnia | 6
compensated respiratory acidosis | 6
electrolyte disturbances | 6
hypomagnesemia | 6
hypophosphatemia | 6
severe hypoalbuminemia | 6
elevated CRP | 6
elevated WBC count | 6
extreme thyroid insufficiency | 6
myxedema | 6
fluid resuscitation | 6
inotropic support | 6
hormonal substitution | 6
intravenous T4 | 6
intravenous T3 | 6
empirical intravenous piperacillin/tazobactam | 6
urine culture | 10
growth of Escherichia coli | 10
material taken from the lower limb wound | 10
growth of Corynobacterium | 10
metronidazole withdrawn | 9
intravenous cefuroxime | 10
intravenous metronidazole | 10
increased CRP level | 16
emergence of clinical and radiological signs of pneumonia | 16
piperacillin/tazobactam | 16
abdomen silent | 16
moderately distended | 16
no signs of bowel movement | 16
enteral nutrition | 16
CT scans of the abdomen | 16
presence of fecal content in the colon and rectum | 16
expansion of the colon and rectum | 16
enhancement and edema of sigmoid and rectal wall | 16
diagnosed bowel obstruction | 16
enemas | 16
violent and abundant diarrhea | 16
inspection of CDI | 16
diagnosis of CDI | 20
PCR test | 20
enteral vancomycin | 20
persistent diarrhea | 24
intravenous metronidazole | 24
enteral fidaxomicin | 24
intravenous tigecycline | 24
piperacillin/tazobactam stopped | 24
no clinical improvement | 31
colonoscopy | 31
extensive swelling of the mucous membrane | 31
no pseudomembranous formations | 31
fecal microbiota transplant | 31
frozen stool from an unrelated healthy donor | 31
donor screened for bacterial pathogens and parasites | 31
transplantation procedure | 31
liquid suspension of donor stool | 31
enema portions | 31
symptoms of diarrhea disappeared | 33
no adverse effects | 33
rapid decrease in CRP levels | 33
recovery from myxedema | 33
discharged to the ordinary ward | 65