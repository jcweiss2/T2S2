78 years old | 0
male | 0
admitted to the hospital | 0
current smoker | 0
hypertension | 0
hyperlipidemia | 0
nifedipine | -2160
candesartan | -2160
atorvastatin | -2160
doxazosin | -2160
sarpogrelate | -2160
levofloxacin eye drops | 0
binocular cataract surgery | 24
fever | 72
dyspnea | 72
cefcapene pivoxil | 72
hypoxia | 72
oliguria | 72
neutrophilia | 72
elevation of the C-reactive protein | 72
impairment of liver and kidney function | 72
bilateral non-segmental consolidation | 72
thickening of the bronchovascular bundles | 72
pleural effusion | 72
tazobactam/piperacillin | 72
continuous hemodiafiltration | 72
ventilatory support | 72
renal function improved | 96
respiratory failure | 96
fever | 96
meropenem | 96
increase in airway pressure | 120
wheezes | 120
corticosteroid treatment | 120
lymphocytes increased | 240
eosinophils increased | 240
nicardipine hydrochloride | 240
sivelestat sodium | 240
levofloxacin injection | 240
respiratory condition worsened | 240
liver dysfunction | 240
steroid therapy | 240
fever continued | 288
levofloxacin eye drops discontinued | 288
fever resolved | 528
respiratory failure resolved | 528
extubated | 528
discharged | 1368
DLST positive | 1368 
drug-induced lung injury | 0