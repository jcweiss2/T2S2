65 years old|0
    male|0
    diabetes|0
    fever|0
    headache|0
    dizziness|0
    cough|0
    fever persists|0
    headache persists|0
    dizziness persists|0
    cough persists|0
    poorly managed diabetes mellitus|-182400
    cranial MRI|0
    multiple abnormal signals|0
    bilateral temporal lobes|0
    hippocampus|0
    sylvian cistern|0
    bilateral cerebellum|0
    fourth ventricle|0
    encephalitis|0
    chest CT scan|0
    multiple lung inflammations|0
    pleural adhesions|0
    pleural effusion|0
    C-reactive protein|0
    CRP 340.0 mg/L|0
    neck stiffness|0
    deep coma|0
    Glasgow Coma Scale score 5|0
    weakness|0
    nausea|0
    repeated vomiting|0
    persistent coma|0
    admission to ICU|0
    lumbar puncture|24
    CSF analysis|24
    CSF cloudiness|24
    CSF white blood cell count 3437/μL|24
    CSF polymorpholeukocytes 85%|24
    CSF glucose 0.6 mmol/L|24
    CSF blood glucose 10.4 mmol/L|24
    CSF microprotein 164.4 mg/dL|24
    Pan's test +++|24
    CSF forceful expulsion|24
    CSF identified as HvKP|48
    virulence factors rmpA|48
    virulence factors iutA|48
    virulence factors iucA|48
    virulence factors iucB|48
    virulence factors iucC|48
    virulence factors iucD|48
    virulence factors iroB|48
    virulence factors iroC|48
    virulence factors iroD|48
    virulence factors fimH|48
    CSF routine|72
    BALF|72
    two sets of blood cultures|72
    HvKP infection|72
    drug sensitivity analysis|72
    resistance to piperacillin|72
    resistance to levofloxacin|72
    sensitivity to amikacin|72
    severe intracranial infection|72
    community-acquired HvKP pathogen|72
    meropenem 2.0 g q8h|72
    intravenous amikacin 0.8 g qd|72
    fever subsided|72
    vital signs stabilized|72
    blood sugar monitoring|72
    blood sugar 6.0–10.0 mmol/L|72
    repeat CSF analysis|216
    CSF clarity|216
    CSF colorlessness|216
    no microorganisms on Gram stain|216
    no CSF culture growth|216
    regained consciousness|264
    endotracheal tube extubated|264
    meropenem treatment 21 days|504
    amikacin treatment 14 days|336
    discharged|288
    