42 years old | 0
female | 0
Systemic Lupus Erythematosus (SLE) | -672
disease modifying drugs | -672
acute calculous cholecystitis | 0
open cholecystectomy | 0
transient leukocytosis | 0
abnormal gall bladder imaging | 0
sepsis | 72
multiorgan dysfunction | 72
catheter-related blood stream infection (CRBSI) | 72
CVC placement in right subclavian vein | -72
CVC removal | 72
new CVC placement in left IJV | 72
free flow of blood from all ports | 72
follow-up chest x-ray normal | 72
correct positioning | 72
absence of pneumothorax | 72
swelling on the left side of neck | 48
local hematoma | 48
catheter removal | 48
new catheter placement in right IJV | 48
dyspnea | 24
desaturation at room air | 24
diminished breath sounds bilaterally | 24
urgent ultrasonography (USG) | 24
chest x-ray | 24
bilateral pleural effusion | 24
pleurocentesis | 24
milky effusion | 24
biochemical analysis | 24
increased triglycerides | 24
bilateral chylothorax | 24
intra pleural drainage tubes placement | 24
under-water seals establishment | 24
chyle drainage | 24
nil per mouth | 24
subjective improvement | 48
total chest tube drainage reduction | 120
drains removal | 216
discharge | 216