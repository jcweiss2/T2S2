41 years old | 0
female | 0
G5P4 | 0
32 weeks pregnant | 0
admitted to the hospital | 0
complaining of dry cough | -72
complaining of shortness of breath | -72
complaining of headache | -72
receiving regular prenatal care | -672
no diabetes mellitus | 0
no hypertension | 0
no bronchial asthma | 0
no other comorbidities | 0
BMI 35.6 | 0
normal blood pressure | 0
heart rate 99 bpm | 0
respiratory rate 24 bpm | 0
oxygen saturations 93-96% | 0
chest x-ray showed diffuse bilateral alveolar infiltrates | 0
diagnosis of sepsis | 0
community acquired pneumonia | 0
started on empiric antibiotic therapy with ceftriaxone | 0
started on empiric antibiotic therapy with azithromycin | 0
COVID-19 PCR swab positive | 0
oxygenation worsened | 15
supplemental oxygen started at 3 L/min | 15
oxygen via high flow nasal cannula started | 24
high flow nasal cannula set at 40 L flow with 100% FiO2 | 24
ABG revealed PaO2 of 111 mmHg | 24
PaO2:FiO2 ratio of 111 | 24
moderate ARDS | 24
transferred to the intensive care unit | 24
repeat ABG revealed PaO2 of 89 mmHg | 31
PaO2:FiO2 ratio of 89 | 31
severe ARDS | 31
dose of furosemide 40 mg given | 31
intravenous dexamethasone started | 31
decision to intubate made | 31
placenta previa with possible accreta | 31
no vaginal bleeding | 31
no signs of fetal distress | 31
endotracheal intubation performed | 35
sevoflurane administered | 35
rocuronium administered | 35
succinylcholine administered | 35
ventilator settings increased to PEEP of 20 cmH2O and FiO2 of 100% | 35
ABG revealed PaO2 of 59 mmHg | 35
PaO2:FiO2 ratio of 59 | 35
sedation initiated with fentanyl and midazolam infusions | 35
repeat ABG revealed PaO2 of 150 mmHg | 37
PaO2:FiO2 ratio of 150 | 37
ventilator settings adjusted | 37
plateau pressure checked and found to be 39 cmH2O | 37
PEEP decreased from 20 cmH2O to 15 cmH2O | 37
vaginal bleeding developed | 38
emergency cesarean section performed | 38
sevoflurane administered | 38
rocuronium administered | 38
midazolam administered | 38
fentanyl administered | 38
oxytocin administered | 38
phenylephrine administered | 38
intravenous bicarbonate administered | 38
baby delivered | 38
baby intubated | 38
Apgar score of 0, 5, and 7 | 38
maternal procedure unremarkable | 38
postoperatively transferred back to the ICU | 38
ventilatory support maintained | 38
ABG performed at 41 hours post-admission | 41
PaO2 of 438 mmHg | 41
PaO2:FiO2 ratio of 438 | 41
plateau pressure 25 cmH2O | 41
convalescent plasma given | 41
oxygenation improved | 65
PEEP and FiO2 weaned down to 10 cmH2O and 40% | 65
ABG demonstrated PaO2 of 92 mmHg | 65
oxygenation continued to improve | 89
ventilator settings gradually weaned | 89
liberated from mechanical ventilation to 3 LPM via nasal cannula | 96
transferred out of the ICU | 96
oxygen requirements continued to improve | 99
transitioned to room air | 99
discharged from the hospital | 288
infant's hospital course notable for negative COVID PCR at 24 and 48 hours post-delivery | 72
infant successfully extubated 48 hours following delivery | 96
placental tissue sent for pathology | 288
placental tissue showed no significant abnormalities | 288