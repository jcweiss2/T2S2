43 years old | 0
female | 0
difficult-to-manage bronchial asthma | -1920
hospitalized | -1920
dry cough | -24
progressive dyspnea | -24
psychomotor agitation | -24
audible wheezing | -24
salbutamol | -24
ipratropium bromide | -24
admitted | 0
diaphoretic | 0
tachycardic | 0
dyspneic | 0
supraclavicular retractions | 0
auscultation with abolished vesicular murmur | 0
Glasgow coma scale 12/15 | 0
arterial blood gases analysis | 0
respiratory acidosis | 0
hypoxemia | 0
invasive ventilatory support | 0
midazolam | 0
propofol | 0
hydrocortisone | 0
magnesium sulfate | 0
antibiotics | 0
cisatracurium | 48
neuromuscular blocking agents | 48
improvement in ABG | 96
ventilatory weaning | 96
dual sedation suspended | 96
NMB suspended | 96
dexmedetomidine | 96
Glasgow coma scale 15/15 | 144
weakness of the neck flexor muscles | 144
facial paresis | 144
muscle strength 1/5 in lower limbs | 144
muscle strength 2/5 in upper limbs | 144
flaccid hyporeflexia | 144
preserved sensitivity | 144
normal cranial nerves | 144
brain MRI | 144
cervical MRI | 144
cerebrospinal fluid study | 144
MRC score 37 points | 144
electromyography | 144
denervation | 144
irritability | 144
polyneuropathic compromise | 144
axonal pattern | 144
ICUAW diagnosis | 144
physiotherapy | 144
comprehensive rehabilitation | 144
ventilator withdrawn | 240
hospital discharge | 720
MRC score 55 points | 720
normal ABG control | 720
symptomatic resolution | 720