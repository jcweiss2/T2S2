61 years old | 0
male | 0
admitted to the hospital | 0
flank pain | -72
dysuria | -72
urgency | -72
frequency | -72
hematuria | -72
fever | -72
chills | -72
rigors | -72
renal colic | -504
nephrolithiasis | -504
staghorn calculus | -504
weight loss | -2160
night sweats | -2160
low grade fevers | -2160
hypotension | 0
hypothermia | 0
urinary tract infection | 0
septic shock | 0
pressor support | 0
norepinephrine | 0
vancomycin | 0
piperacillin-tazobactam | 0
ill-defined liver lesions | 0
liver biopsy | 216
bone marrow biopsy | 216
Hodgkin lymphoma | 216
chemotherapy | 216
doxorubicin | 216
dacarbazine | 216
vinblastine | 216
bleomycin | 216
shortness of breath | 120
hypoxia | 120
fluid overload | 120
lasix | 120
colonoscopy | 144
esophago-gastro-duo-denoscopy | 144
tubular adenoma | 144
gastric folds | 144
chronic gastritis | 144
discharged | 216
readmitted | 264
fever | 264
weakness | 264
fatigue | 264
liver enzymes | 0
alkaline phosphatase | 0
alanine transaminase | 0
aspartate transaminase | 0
total protein | 0
albumin | 0
urine dipstick | 0
urine microscopy | 0
cortisol level | 0
TSH | 0
Free T4 | 0
blood culture | 0
urine culture | 0
CT scan | 0
trans-thoracic echocardiogram | 120
Reed-Sternberg cells | 216
CD15 | 216
CD30 | 216
CD45 | 216
CD3 | 216
CD20 | 216
immunohistochemical stains | 216
staging | 216
CT Chest | 216
hilar lymphadenopathy | 216
pulmonary function test | 216
smoking | -10080
alcohol consumption | -10080
nephrolithiasis | -10080
lithotripsy | -10080
family history | 0
medication history | 0
HIV ELISA | 0
sedimentation rate | 0
C-Reactive Protein | 0
hepatitis B | 0
hepatitis A | 0
hepatitis C | 0
ANA panel | 0
ANCA panel | 0
rheumatoid factor | 0
C3 | 0
C4 | 0