38 years old | 0
    male | 0
    Hepatitis B Virus (HBV) infection | -4320
    Polyarteritis Nodosa (PAN) | -4320
    weight loss | -8760
    myalgias | -8760
    fever | -8760
    skin erythema | -8760
    deterioration of renal function | -8760
    new onset of diabetes mellitus Type II | -8760
    hypertension | -8760
    chronic renal failure | -4320
    diabetes mellitus Type II | -4320
    prednisolone | -4320
    cyclophosphamide | -4320
    Tenofovir | -4320
    discontinued Tenofovir | -2016
    acute abdomen | 0
    septic shock | 0
    free sub diaphragmatic air | 0
    laparotomy | 0
    peritonitis | 0
    three perforations of the small intestine | 0
    segmental enterectomy | 0
    anastomosis | 0
    mechanical ventilation | 0
    circulatory support | 0
    acute-on-chronic renal failure | 0
    weaned off ventilator | 72
    haemodynamically stable | 72
    started Tenofovir | 168
    IV methylprednisolone | 168
    abdominal drain catheter presented enteric content | 168
    second explorative laparotomy | 168
    two new perforations | 168
    multiple areas of patchy necrosis | 168
    suture repair | 168
    open abdomen | 168
    vacuum device | 168
    plan for re-laparotomy | 168
    plasma exchanges | 168
    IV cyclophosphamide | 168
    IV methylprednisolone | 168
    IV prednisone | 168
    third laparotomy | 216
    three new necrotic lesions | 216
    suture repair | 216
    necrotic lesion on left lobe of liver | 216
    fourth laparotomy | 264
    segmental enterectomy | 264
    anastomosis | 264
    cholecystectomy | 264
    anastomotic leak | 264
    gangrenous gallbladder | 264
    died | 360
    septic shock | 360
    multiple organ failure | 360