74 years old| 0
man | 0
presented to the emergency department | 0
diarrhoea | -72
vomiting | -72
pansystolic murmur | 0
Janeway lesion | 0
Osler node | 0
nail bed haemorrhage | 0
amalgam restoration | 0
absent upper first premolar | 0
absent upper left molar | 0
elevated inflammatory markers | 0
Staphylococcus aureus bacteraemia | 0
severe mitral regurgitation | 0
vegetations on mitral valve | 0
vegetations on aortic valve | 0
renal failure | 0
worsening sepsis | 0
anuric | 192
haemodialysis | 192
haemodialysis | 216
transferred to tertiary hospital | 240
admitted to intensive care unit | 240
continuous venovenous haemofiltration | 240
positive SARS-CoV-2 nasopharyngeal swab | 264
nausea | 576
vomiting | 576
peripheral ground glass change | 576
bilateral pleural effusions | 576
COVID-19 pneumonia | 576
supplementary oxygen | 576
oral dexamethasone | 576
intravenous remdesivir | 576
acute respiratory distress syndrome | 744
death | 744
- 74 years old | 0
7 man | 0
renal failure | 120
worsening sepsis | 120
- male | 0
- presented to the emergency department | 0
- diarrhoea | -72
. vomiting | -72
- agitated | 0
$ GCS 12/15 | 0
- pansystolic murmur | 0
- Janeway lesion | 0
0 Osler node | 0
- nail bed haemorrhage | 0
- amalgam restoration | 0
- absent upper first premolar | 0
- absent upper left molar | 0
- elevated inflammatory markers | 0
- blood cultures taken | 0
- started on intravenous ceftriaxone | 0
(blood culture grew Staphylococcus aureus | 0)
- severe mitral regurgitation | 0
8 vegetations on mitral valve | 0
- vegetations on aortic valve | 0
- negative SARS-CoV-2 swab | 0
- renal failure | 120
- worsening sepsis | 120
- anuric | 192
- haemodialysis | 192
- haemodialysis | 216
- transferred to tertiary hospital | 240
# admitted to intensive care unit | 240
- continuous venovenous haemofiltration | 240
- positive SARS-CoV-2 swab | 264
- nausea | 576
- vomiting | 576
- peripheral ground glass change | 576
- bilateral pleural effusions | 576
- COVID-19 pneumonia | 576
! supplementary oxygen | 576
- oral dexamethasone | 576
- intravenous remdesivir | 576
- acute respiratory distress syndrome | 744
- death | 744
