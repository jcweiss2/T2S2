43 years old | 0
male | 0
Caucasian | 0
admitted to the Emergency Department | 0
fever | -48
sneezing | -48
fatigue | -48
sore throat | -48
dry cough | -48
no dyspnea | -48
mild cognitive impairment | -6480
arterial hypertension | -6480
systemic lupus erythematosus | -4896
lupus nephritis | -4896
mycophenolate | -4896
prednisone | -4896
family history negative for cancer | 0
family history negative for endocrinopathy | 0
family history negative for inflammatory diseases | 0
parents dead | 0
no children | 0
physical examination on admission | 0
fever (38 °C) | 0
oxygen saturation of 94% | 0
respiratory rate of 18 breaths/min | 0
decreased breath sounds | 0
coarse crackles in both lung bases | 0
white blood cell count of 7110/μL | 0
mild lymphocytopenia 650/μL | 0
D-dimer 0.73 μg/ml | 0
C-reactive protein 62 mg/L | 0
PCT 94 ng/mL | 0
hemoglobin normal | 0
platelets normal | 0
serum electrolytes normal | 0
creatinine normal | 0
liver function test normal | 0
arterial blood gas analysis | 0
pH 7.44 | 0
pO2 75 mm Hg | 0
pCO2 37 mm Hg | 0
SARS-Cov-2 RNA positive | 0
chest computed tomography scan | 0
bilateral ground-glass opacities | 0
hyperdense and irregular foci in the thoracic vertebral bodies | 0
empirical antibiotic therapy with piperacillin/tazobactam | 0
oxygen support | 0
general condition improved | 288
C-reactive protein normalized | 288
blood and urine culture tests negative | 288
PCT remained elevated (84 ng/mL) | 288
serum CTN measured | 288
CTN 2120 pg/mL | 288
carcinoembryonic antigen 108 ng/mL | 288
total and ionized calcium normal | 288
thyrotropin normal | 288
thyroxine normal | 288
neck examination | 288
painless right laterocervical swelling | 288
neck ultrasound | 288
inhomogeneously echogenic lymph nodes | 288
small punctate calcifications | 288
nonhomogeneous thyroid | 288
multiple nodules | 288
cytologic examination by fine-needle aspiration | 288
MTC diagnosis | 288
CTN value in the aspiration needle washout fluid >2000 pg/mL | 288
PCT:CTN ratio 3.96 | 288
neck, lung, and abdomen computed tomography scan | 288
no lesions other than in the neck lymph nodes | 288
multiple sclerotic lesions at dorsal spine level | 288
multiple sclerotic lesions at hip bone level | 288
fluorine-18 fluorodeoxyglucose positron emission tomography/computed tomography scan | 288
increased tracer uptake in the right laterocervical lymph nodes | 288
total thyroidectomy with bilateral cervical lymph node dissection | 432
histologic examination of the surgical specimen | 432
MTC confirmed | 432
neoplastic cells positive for CTN, carcinoembryonic antigen, synaptophysin, chromogranin A, and thyroglobulin | 432
MTC metastases in 3 of 12 lymph nodes | 432
pathologic T1b-N1a, stage III | 432
blood tests 48 hours after surgery | 480
CTN 986 pg/mL | 480
PCT 16 ng/mL | 480
nasopharyngeal and oropharyngeal swabs negative | 528
discharged | 528
oral therapy of prednisone | 528
oral therapy of ramipril | 528
oral therapy of levothyroxine | 528
oral therapy of cholecalciferol | 528
oral therapy of calcium carbonate | 528
6-month follow-up | 4320
(18)F-fluorodihydroxyphenylalanine positron emission tomography | 4320
no suspicious fixations at the thyroid lodge and cervical lymph node stations | 4320
multiple osteoblastic foci in the skeletal area | 4320
CTN 921 pg/mL | 4320
PCT 16 ng/mL | 4320
close follow-up planned | 4320