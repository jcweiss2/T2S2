32 years old | 0
female | 0
34 weeks of gestation | 0
admitted to the ICU | 0
severe coronavirus disease 2019 | 0
hypoxemic respiratory failure | 0
SpO2: 94% | 0
oxygen therapy by reservoir bag at 15 L/min | 0
respiratory rate of 30 breaths per min | 0
piperacillin–tazobactam | 0
methylprednisolone | 0
remdesivir | 0
high-flow nasal cannula therapy | 0
intubated | 6
persistent hypoxemic respiratory failure | 6
standard lung-protective ventilation | 6
pregnancy terminated | 6
acute respiratory distress syndrome | 6
fetal distress | 6
lower segment cesarean section | 6
live female baby delivered | 6
PaO2/FiO2 ratio post LSCS was 120 | 6
prone ventilation sessions | 6
diffuse subcutaneous edema of the face | 12
subcutaneous edema reduced | 16
percutaneous tracheostomy | 168
septic shock with Klebsiella pneumoniae bacteremia | 168
antimicrobials | 168
colistin | 168
meropenem | 168
shock recovered | 336
weaning initiated | 384
spontaneous breathing trial | 384
inability to close left eyelid | 384
deviation of the angle of mouth to the right side | 384
no other focal neurological deficit | 384
plantar reflexes were of flexor response | 384
examination of both ears did not reveal any discharge | 384
power of all four limbs was reduced | 384
Medical Research Council sum score of 40 | 384
diagnosis of critical illness neuromyopathy | 384
patching of the eyelid | 384
lubrication with eye drops | 384
contrast-enhanced computed tomography scan | 384
soft-tissue swelling with fat stranding in the left cheek and masseter muscle | 384
no evidence of stroke | 384
no significant compression in the tract of the facial nerve | 384
no fracture or any osseous lesion in the facial canal | 384
active limb physiotherapy | 384
good glycemic control | 384
steroids deferred | 384
acyclovir not administered | 384
improvement in neuromuscular strength | 552
weaned from mechanical ventilation | 552
decannulated | 720
left facial nerve palsy persisted | 720
House–Brackmann Facial Nerve Grade IV | 720
magnetic resonance imaging of the brain with contrast | 720
subtle postcontrast enhancement in the cisternal and intracanalicular part of the 7th and 8th nerve complex | 720
discharged home | 720
complete resolution of paresis | 1440
no serious long-term effects like crocodile tears syndrome | 1440