52 years old | 0
male | 0
admitted to the hospital | 0
body mass index 23.6 kg/m2 | 0
no comorbidities | 0
open modified Scopinaro procedure | -7200
weight 216 kg | -7200
BMI 57.4 kg/m2 | -7200
weight reganance | -2400
incisional hernia | -2400
bariatric revisional surgery | -2400
hernia repair | -2400
weight 170 kg | -2400
BMI 45.1 | -2400
gastric pouch leak | -2400
intra-abdominal collections | -2400
sepsis | -2400
conservative management | -2400
open abdomen | -2400
negative wound pressure therapy | -2400
parenteral nutrition | -2400
intravenous antibiotics | -2400
epithelized gastrocutaneous fistula | -1200
controlled but persistent drainage | -1200
proximal edge of planned ventral hernia | -1200
upper endoscopy | -1200
fistulous orifice | -1200
vertical staple line | -1200
esophagogastric junction | -1200
extraluminal extravasation | -1200
recurrent left subphrenic abscess | -1200
endoscopic treatment | -1200
argon plasma coagulation | -1200
internal drainage | -1200
external drainage | -1200
clipping | -1200
fibrin sealants | -1200
e-vac therapy | -1200
stenting | -1200
multidisciplinary team discussion | 0
decision to proceed with innovative endoscopic technique | 0
placement of CSDO | 0
Occlutech muscular VSD occluder | 0
intravenous sedation | 0
topic anesthesia | 0
fistula cannulation | 0
biliary stent deployment system | 0
direct endoscopic guidance | 0
extraluminal leakage | 0
contrast injection | 0
Amplatz extra stiff guidewire | 0
fluoroscopy | 0
delivery system | 0
CSDO deployment | 0
endoscopic guidance | 0
fluoroscopic guidance | 0
no immediate adverse events | 0
contrast study | 0
no extravasation of contrast material | 0
restricted oral intake | 24
liquid diet | 24
regular diet | 288
pigtail drain | 0
accidental displacement of pigtail | 432
systemic signs of sepsis | 432
computed tomography | 432
fluoroscopy | 432
recurrence of abscess | 432
partial dislodgment of CSDO | 432
second attempt with oversized disc | 432
Occlutech Figulla Flex II UNI | 432
sealing of fistulous orifice | 432
upper endoscopy | 1296
contrast-enhanced CT scan | 1296
device engrafted | 1296
reduction of chronic abscess | 1296
no signs of fistula recurrence | 1296
pigtail removal | 1296
no drainage | 1296