77 years old | 0
male | 0
admitted to ICU | 0
confusion | 0
shortness of breath | 0
tachycardia | 0
hypothermia | 0
hypotension | 0
pre-diagnosis of acute respiratory failure | 0
pre-diagnosis of SIRS | 0
intubated | 0
connected to ventilator | 0
decrease in respiratory sounds | 0
coarse rales | 0
prolongation of expirium | 0
bilateral biphasic expiratory ronchi | 0
obstructive pattern on pulmonary function test | -120
history of tuberculosis | -8760
history of COPD | -8760
history of Hyperthyroidism | -8760
history of Diabetes Mellitus | -8760
Glasgow Coma Score 6 | 0
APACHE II 34 | 0
MODS 8 | 0
pulse 122/min | 0
arterial blood pressure 82/41 mmHg | 0
respiratory rate 30/min | 0
temperature 35°C | 0
Leukocyte 27600/mm3 | 0
C-reactive protein 52 mg/L | 0
thyrotoxicosis | 0
free thyroxine 8.5 ng/dL | 0
thyrotropin < 0.05 μIU/mL | 0
thyroid receptor antibodies 0.9 IU/mL | 0
thyroid ultrasonography showed solid hyperechoic nodule | 0
treatment with propranolol | 0
treatment with methimazole | 0
pneumonic infiltration on chest X-ray | 0
increase in ground glass density on chest X-ray | 0
no pathology on ECG | 0
diastolic dysfunction on Echocardiography | 0
fever 38.4°C | 48
Ampicilline-Sulbactam treatment | 48
Levofloxacin treatment | 48
no growth on cultures | 48
substituted treatment with Piperacilline/Tazobactam | 168
substituted treatment with Trimetoprim/Sulfametaxazol | 168
substituted treatment with Claritromycin | 168
bronchoscopy | 168
fungus ball seen on thoracic CT | 168
narrow lumens of trachea and bronchi | 168
diffuse white-colored plaques | 168
thin-walled necrotic lesion on thorax CT | 168
crescent sign on thorax CT | 168
histopathological examination showed mixed active inflammation | 168
histopathological examination showed fibrous scarring | 168
histopathological examination showed microscopic abscess cavity | 168
histopathological examination showed central bronchiectasis | 168
histopathological examination showed dense peribronchial inflammation | 168
histopathological examination showed fungus ball | 168
histopathological examination showed septate hyphae of Aspergillus fumigatus | 168
Aspergillus fumigatus grew on BAL culture | 168
voriconazole treatment | 168
loading dose of voriconazole 1×400 mg i.v. | 168
maintenance dose of voriconazole 2×200 mg i.v. | 168
disease became more severe | 432
multiple organ failure | 432
death | 432