56 years old | 0
female | 0
admitted to the hospital | 0
weakness | -720
numbness | -720
lower extremities weakness | -720
hands weakness | -720
neck weakness | -720
type 2 diabetes mellitus | 0
hypertension | 0
necrotizing pancreatitis | -8760
gallstones | -8760
total parenteral nutrition (TPN) | -2190
discontinued TPN | -168
normal diet | -168
Guillain-Barré syndrome (GBS) | -720
albuminocytologic dissociation | 0
lumbar puncture | 0
brain magnetic resonance imaging (MRI) | 0
small vessel ischemic changes | 0
intravenous immunoglobulin (IVIG) treatment | 0
encephalopathy | 120
pancytopenia | 120
hypotensive | 120
blood pressure 64/48 mmHg | 120
unresponsive to verbal stimuli | 120
minimally responsive to painful stimuli | 120
Glasgow Coma Scale (GCS) score of 6 | 120
anasarcic | 120
flaccid paralysis | 120
malnourished | 120
septic state | 120
calcium 6.7 mg/dL | 120
hemoglobin 9.4 g/dL | 120
white cell count 2.1×10^9/L | 120
phosphorus 1.1 mg/dL | 120
creatinine <0.2 mg/dL | 120
albumin <1.5 gm/dL | 120
lactate 4 mmol/L | 120
Nutritional risk screening (NRS-2002) score of 5 | 120
malnutrition universal screening (MUST) score of 5 | 120
intubated | 120
intravenous fluids | 120
norepinephrine | 120
meropenem | 120
vancomycin | 120
anidulafungin | 120
sepsis | 120
empirical treatment with high-dose intravenous thiamine | 120
electroencephalogram (EEG) | 168
diffuse slow waves | 168
severe metabolic encephalopathy | 168
brain MRI | 216
hyperintensity of the bilateral medial thalamus | 216
Wernicke’s encephalopathy | 216
serum thiamine level 104 nmol/L | 216
improved mental status | 288
able to understand simple commands | 288
discontinued norepinephrine | 288
discontinued antimicrobial treatment | 288
extubated | 360
electromyography (EMG) | 504
severe sensorimotor polyneuropathy | 504
transferred out of the intensive care unit (ICU) | 1008
thiamine supplementation continued | 1008
dry beriberi | 0
ascending neuropathy | 0
paralysis | 0
Wernicke’s encephalopathy | 0
thiamine deficiency | 0
malabsorption | 0
alcohol abuse | 0
anorexia nervosa | 0
dieting | 0
bariatric surgery | 0
diarrhea | 0
celiac disease | 0
tropical sprue | 0
dysentery | 0
burns | 0
pregnancy | 0
dialysis | 0
malignancy | 0
cardiomyopathy | 0
cardiomegaly | 0
heart failure | 0
dyspnea | 0
peripheral edema | 0
Shoshin beriberi | 0
cardiogenic shock | 0
lactic acidosis | 0
multi-organ failure | 0
ataxia | 0
ophthalmoplegia | 0
nystagmus | 0
irreversible cognitive impairment | 0
magnetic resonance imaging (MRI) | 0
serum thiamine levels | 0
axonal abnormalities | 0
impaired acetylcholine transmission | 0
axonal injuries | 0
painful sensory or sensorimotor polyneuropathy | 0
muscle weakness | 0
Guillain-Barré syndrome (GBS) | 0
acute inflammatory demyelinating polyradiculoneuropathy (AIDP) | 0
infection | 0
electromyography | 0
albuminocytologic dissociation | 0
cerebrospinal fluid | 0
white blood cells | 0
chronic inflammatory demyelinating polyneuropathy (CIDP) | 0
cranial nerves | 0
bulbar nerves | 0
autonomic instability | 0
critical illness myopathy | 0
critical illness polyneuropathy | 0
sepsis | 0
encephalopathy | 0
delirium | 0
mechanical ventilation | 0
neuromuscular impairment | 0
cognitive impairment | 0
thiamine supplementation | 0
high-dose thiamine | 0
magnetic resonance imaging (MRI) | 0
electrophysiological studies | 0
alcohol abuse | 0
severe protein-calorie malnutrition | 0
bariatric surgery | 0
total parenteral nutrition (TPN) | 0
malabsorption | 0
increased caloric requirements | 0
neuropathy | 0
weakness | 0
cardiomyopathy | 0
autonomic instability | 0