66 years old | 0
female | 0
admitted to hospital | 0
lower abdominal pain | -24
vital signs within normal range | -24
urine/blood investigations unremarkable | -24
CT abdomen/pelvis | -24
large right sided pelvi-ureteric junction calculus | -24
xanthogranulomatous pyelonephritic kidney | -24
elective surgery planned | -24
endoscopic procedure consented | -24
ureteropyeloscopy and lasertripsy surgery | -72
mixed growth in urine culture | -72
polyps in right ureter | -72
pus in renal pelvis | -72
intraoperative retrograde pyelogram | -72
no evidence of fistula | -72
ureteric stent inserted | -72
discharged with oral antibiotics | -72
ureteric biopsies showed inflammatory changes | -72
repeat pyeloscopy procedure | -120
renal calculi treated with lasertripsy | -120
ureteric stent inserted | -120
intraoperative RPG unremarkable | -120
ureteric stent removed | -113
severe sepsis | 0
hypothermia | 0
hypotension | 0
tachycardia | 0
tachypnoea | 0
elevated inflammatory markers | 0
moderate renal impairment | 0
positive urinalysis | 0
leukocytes in urine | 0
nitrites in urine | 0
blood in urine | 0
urine culture showed mixed growth | 0
blood cultures showed Proteus mirabilis | 0
CT KUB showed peri-nephric stranding | 0
emergency cystoscopy | 0
RPG showed uretero-duodenal fistula | 0
stent insertion | 0
transfer to intensive care unit | 0
right sided nephrectomy | 24
laparoscopic approach | 24
conversion to open surgery | 24
adhesiolysis and haemostasis | 24
no resection of duodenum | 24
post-operative management | 24
tolerating fluids on Day 3 | 72
full diet on Day 5 | 120
discharged home | 168
follow-up appointment | 4320
no urinary symptoms | 4320
no pain issues | 4320
CT abdomen/pelvis showed no abnormal collections | 4320