72 years old | 0
male | 0
admitted to the hospital | 0
fever | -12
chills | -12
cough | -12
chest pain | -12
total leucocyte count 37 100/mm3 | -12
consolidation in the right lung | -12
low blood pressure | -12
noradrenaline infusion started | 0
peripherally placed 18G intravenous cannula | 0
broad-spectrum antibiotics | 0
fluid resuscitation | 0
vasopressor support | 0
blood pressure stabilized | 2
vasopressor tapered off | 2
CVC placement not attempted | 2
swelling over the dorsum of the left hand | 12
purplish discoloration | 12
infusion stopped | 12
IV cannula removed | 12
new IV cannula placed | 12
NA infusion tapered off | 16
NA infusion stopped | 16
topical nitroglycerin applied | 12
topical nitroglycerin repeated | 16
hand elevated | 12
heat application | 12
swelling and discoloration improved | 48
skin texture near normal | 48
phentolamine not available | 0
terbutaline not available | 0
discharged | 60