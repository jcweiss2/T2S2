57 years old | 0
male | 0
admitted to the hospital | 0
breathlessness | -96
abdominal discomfort | -96
40-pack year smoking history | 0
febrile | 0
tachycardic | 0
lactate 4 mmol/l | 0
colonoscopy | -120
biopsy of a splenic flexure polyp | -120
diverticular disease | -120
diagnosis of possible abdominal perforation and sepsis | 0
deteriorated | 24
painful cold legs | 24
hypotensive | 24
agitated | 24
sweaty | 24
peripheral mottling | 24
massive hepatomegaly | 24
lactate 14 mmol/l | 24
hypoglycaemia | 24
resuscitated with crystalloid and dextrose | 24
transferred to the ICU | 24
cardiac arrest | 24
pulseless electrical activity | 24
intubated | 24
cardiopulmonary resuscitation | 24
return of spontaneous circulation | 24
central venous catheter inserted | 24
right internal jugular vein large and non-compressible | 24
central venous pressure 31 mmHg | 24
consumptive coagulopathy | 24
INR 5.9 | 24
fibrinogen 0.2 g/l | 24
platelets 38×10^9/l | 24
transthoracic echo | 24
massive pericardial effusion | 24
right ventricular collapse | 24
electrocardiogram | 0
electrical alternans | 0
chest X-ray | 0
enlarged heart shadow | 0
pericardial effusion drained | 24
700 ml of fluid aspirated | 24
pericardial fluid heavily blood stained | 24
cytological examination not possible | 24
CT of the chest, abdomen and pelvis | 48
CT aortogram | 48
haematoma in the distal arch of the aorta | 48
haematoma in the descending aorta | 48
type A dissection not excluded | 48
transoesophageal echocardiogram | 60
type A dissection excluded | 60
dissection flap in the descending aorta | 60
left-sided pleural effusion | 60
colour flow Doppler | 60
true lumen | 60
cardiovascular support | 72
respiratory support | 72
renal support | 72
serial echocardiograms | 72
moderate recurrence of the pericardial effusion | 72
no significant haemodynamic compromise | 72
paraplegia | 168
pleural effusion | 168
pleural effusion drained | 168
pleural fluid showed cells with positive epithelial and mesothelial immunostains | 168
metastatic adenocarcinoma | 168
primary lung tumour | 168
suspicious spiculate lesion in the left upper lobe | 168
died | 1440
lung cancer | 0 
symptomatic pericardial effusion | 0 
type B aortic dissection | 0