35 years old | 0
female | 0
scheduled for resection of giant cell tumor | 0
resection of giant cell tumor of the right hand radius bone | 0
arthroplasty | 0
coagulation profile were within the normal limits | -24
preoperative routine investigations were within the normal limits | -24
monitored for heart rate | 0
monitored for electrocardiography | 0
monitored for noninvasive blood pressure | 0
monitored for pulse oximetry | 0
peripheral intravenous access was secured | 0
right supraclavicular brachial plexus block was performed | 0
paresthesia technique using anatomical landmarks | 0
combination of 0.5% bupivacaine and 2% lignocaine with adrenaline | 0
complained of slight chest pain | 0
chest expansion and air entry was bilaterally equal | 0
X-ray chest performed showed no pneumothorax or fluid collection | 0
sedated with 1 mg of injection midazolam | 0
surgery was allowed to commence | 0
surgery lasted about one and half hours | 1.5
patient was shifted to the recovery room | 1.5
patient remained symptom free except for slight chest discomfort | 1.5
vitals were stable | 1.5
ECG showed normal sinus rhythm | 1.5
repeat supine X-ray chest was again insignificant | 1.5
supplemented with oxygen | 1.5
adequate sedation and analgesia was ensured | 1.5
shifted from postanesthesia care unit to her ward | 1.5
patient remained symptom free for another 12–14 h | 12
started complaining chest pain and palpitation | 12
increasing severity of chest pain and palpitation | 12
significant reduction in chest expansion on the right side | 12
air entry was almost absent on the right side | 12
X-ray chest showed a massive fluid collection on the right side | 12
partial collapse of the right lung | 12
shifted to operation theater | 12
intercostal tube drainage was inserted | 12
approximately 1300 ml of collected blood was drained out | 12
blood samples were sent for cross matching | 12
emergency investigations were sent | 12
arterial gas analysis showed a mixed picture | 12
compensated metabolic acidosis with respiratory alkalosis | 12
evacuation of hemothorax | 12
patient symptoms improved significantly | 12
administered 4 units of fresh whole blood | 12
shifted to intensive care unit | 12
nursed in propped up position | 12
oxygen was given | 12
analgesic was given | 12
antibiotics cover was given | 12
stable vitals after stay of 5 days in ICU | 60
X-ray chest revealed almost complete expansion of the right lung | 60
retained part of hemothorax | 60
CT guided thoracoscopic evacuation | 60
discharged on tenth postoperative day | 120
satisfactory condition | 120