25 years old | 0
female | 0
Hispanic | 0
sacral myofibroblastic sarcoma | -672
sacrectomy | -672
lumbopelvic fixation | -672
hardware revisions | -336
iliac screw revision | -336
intrathecal pain pump placement | -336
neck pain | 0
headache | 0
fever | 0
somnolent | 0
seizure | 0
lorazepam | 0
levetiracetam | 0
nonspecific hypodensities | 0
lumbar puncture | 0
broad-spectrum antibiotics | 0
intubated | 0
depressed level of consciousness | 0
electroencephalogram | 0
mild generalized slowing | 0
left temporal dysfunction | 0
no epileptiform discharges | 0
cerebrospinal fluid examination | 0
WBC count 5781 mm3 | 0
protein 578 mg/dL | 0
glucose <30 mg/dL | 0
Gram-negative rods | 0
E. coli | 0
K1 strain | 0
intrathecal pump removal | 24
wound culture | 24
E. coli | 24
Candida parapsilosis | 24
fluconazole | 24
MRI brain | 24
multifocal bilateral cerebral and cerebellar cortically based nonenhancing diffusion restricting lesions | 24
cortical infarcts | 24
microhemorrhage | 24
no leptomeningeal enhancement | 24
CT angiogram | 48
no arterial occlusion | 48
no stenosis | 48
no dissection | 48
no vasospasm | 48
transthoracic echocardiogram | 48
unremarkable | 48
transesophageal echocardiogram | 48
not pursued | 48
MRI brain venogram | 48
no dural venous sinus thrombosis | 48
extubated | 96
mild encephalopathy | 96
no focal findings | 96
meropenem | 0
ceftriaxone | 96
meningeal doses | 96
cefepime | 96
hardware infection | 96
discharged | 384
phenytoin | 384
ceftriaxone | 384
cefepime | 384
phenytoin stopped | 408
good recovery | 408
no neurological deficits | 408