28 years old | 0
female | 0
referred to hospital | -3024
singleton pregnancy | -3024
conceived through IVF-ET | -3024
sudden uterine contraction | -720
genital bleeding | -720
watery discharge | -720
speculum examination | -720
positive monoclonal antibodies against insulin-like growth factor-binding protein 1 | -720
suspected premature rupture of the membrane | -720
temperature over 38°C | -720
tachycardia | -720
uterine tenderness | -720
intravenous ampicillin | -720
gentamicin | -720
amniocentesis | -720
blood culture | -720
vaginal discharge culture | -720
early premature rupture of the membrane | -720
blue-green vaginal discharge | -720
indigo carmine injection | -720
elevated white blood cell count | -720
elevated C-reactive protein level | -720
amniotic fluid inflammatory cells | -720
Candida glabrata in amniotic fluid | -720
Candida glabrata in vaginal discharge | -720
temperature over 38°C persisted | -720
1,3:β-D-glucan negative | 0
candidemia not suspected | 0
decision to terminate pregnancy | 24
delivery | 24
fever resolved | 24
Candida glabrata in blood culture | 192
readmission | 192
absence of fever | 192
uterine tenderness | 192
elevated inflammatory markers | 192
systemic candidiasis | 192
candida endophthalmitis | 192
intravenous fluconazole | 192
chorioamnionitis confirmed by histology | 192
maternal inflammatory response stage II grade I | 192
fetal inflammatory response stage I grade I | 192
Candida spp. in chorion | 192
neutrophilic infiltration in chorion | 192
