62 years old | 0
    male | 0
    penetrating trauma in right chest | 0
    left pneumonectomy due to pulmonary tuberculosis infection | -209952
    pulmonary tuberculosis infection | -209952
    symptoms of dyspnea | -72
    symptoms of hemoptysis | -72
    respiratory rate 23 breaths per minute | 0
    oxygen saturation 90% in room air | 0
    conscious | 0
    fully responsive to questions | 0
    initial vital signs stable | 0
    blood pressure 150/90 mm Hg | 0
    heart rate 100 beats per minute | 0
    no use of inotropic drugs | 0
    hemoglobin level 12.2 g/dL | 0
    partial oxygen pressure 60 mm Hg | 0
    chest computed tomography | 0
    foreign body in medial basal segment of right lower lobe | 0
    fracture of right seventh rib | 0
    no pneumothorax | 0
    no hemothorax | 0
    dyspnea ongoing | 0
    hemoptysis ongoing | 0
    foreign body could cause additional lung parenchymal damage | 0
    foreign body could cause infection | 0
    decided to perform emergent surgery | 0
    general anesthesia | 0
    intermittent apnea technique | 0
    mini-thoracotomy via right mid-axillary line of sixth intercostal space | 0
    adhesiolysis of whole lung field | 0
    retracted lung toward apex | 0
    identified opening site of penetration tract at right lower lobe medial basal segment | 0
    no damage to major vessels | 0
    no damage to hilar structure airways | 0
    Duval clamps placed parallel to wound tract | 0
    linear stapler placed through tract | 0
    fired stapler to separate lung parenchyma | 0
    exposed bleeding focus | 0
    exposed injured airway | 0
    hemostasis achieved with multiple 3-0 polypropylene interrupted-suture ligation | 0
    airway control achieved with multiple 3-0 polypropylene interrupted-suture ligation |'0
    extracted 1.3-cm metal fragment at end of distal wound tract | 0
    indwelled 28-Fr right-angled chest tube in right pleural cavity | 0
    wound closed in standard manner | 0
    total surgery time 90 minutes | 0
    no transfusion during surgery | 0
    endotracheal tube removed | 0
    transferred to general ward | 0
    recovered from general anesthesia | 0
    no significant complications after surgery | 0
    chest tube removed on third day of admission | 72
    discharged on seventh day of admission | 168
    no notable events after surgery | 168
    no additional transfusions | 168

