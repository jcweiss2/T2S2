65 years old | 0
woman | 0
scheduled to undergo a left lobe hepatectomy | 0
hepatocellular carcinoma | 0
liver cirrhosis | 0
Child-Pugh class A | 0
chronic hepatitis B | 0
intravenous glycoppyrolate 0.2 mg | -240
general anesthesia induced | -240
propofol 100 mg | -240
rocuronium 50 mg | -240
remifentanil 40 µg | -240
sevoflurane 1-2.5% | -240
remifentanil 0.1-0.25 µg/kg/min | -240
rocuronium 5-10 µg/kg/min | -240
intubated | -240
ventilated mechanically | -240
monitored by EKG | -240
arterial blood pressure | -240
central venous pressure | -240
SpO2 | -240
vital signs stable | -240
hepatectomy with CUSA® started | -1
sudden decrease in arterial blood pressure | 0
systolic blood pressure <40 mmHg | 0
end-tidal carbon dioxide <26 mmHg | 0
SpO2 <50% | 0
tachycardia 1100-135 beats/min | 0
ST elevation on EKG | 0
resuscitation with colloid | 0
catecholamines administration | 0
intravenous epinephrine 1 mg | 0
norepinephrine infusion | 0
intraoperative ultrasonography revealed air emboli | 0
diagnosed with VAE | 0
diagnosed with PAE | 0
arterial blood gas analysis at diagnosis | 0
pH 7.278 | 0
pCO2 51.3 mmHg | 0
PO2 84.6 mmHg | 0
HCO3- 24.2 mmHg | 0
SaO2 94.4% | 0
FiO2 0.5 | 0
systolic blood pressure maintained at 90 mmHg | 10
heart rate maintained at 110 beats/min | 10
central venous pressure 2 mmHg | 10
end-tidal carbon dioxide restored to 32 mmHg | 10
ABGA at 30 minutes after episode | 30
pH 7.338 | 30
pCO2 44.3 mmHg | 30
PO2 234.0 mmHg | 30
HCO3- 24.0 mmHg | 30
SaO2 99.6% | 30
FiO2 1.0 | 30
norepinephrine infusion continued | 70
fluid resuscitation continued | 70
colloid 1000 ml | 70
crystalloid 500 ml | 70
air emboli in left heart disappeared | 70
attempt to aspirate air with jugular catheter | 70
hepatectomy restarted | 70
hepatectomy completed | 70
systolic pressure maintained at 90 mmHg | 70
total anesthesia time 5 hours | 300
total fluid administered 2950 ml | 300
total urinary output 220 ml | 300
total blood loss 800 ml | 300
postoperative intubation | 300
postoperative mechanical ventilation | 300
response only to intense pain | 300
systolic pressure maintained at 90 mmHg | 300
postoperative PT/PTT 25.5/51.8 sec | 300
fibrinogen 96 mg/dl | 300
d-dimer 6519 ng/ml | 300
antithrombin III 19% | 300
CK-MB 40.74 ng/ml | 300
troponin-T 1.880 ng/ml | 300
postoperative EKG ST elevation in II, III, aVF | 300
POD 1 EKG normal | 24
trans-thoracic echocardiogram unremarkable | 24
no PFO identified | 24
vital signs stable | 24
norepinephrine tapered out | 24
POD 5 mental status unchanged | 120
brain CT multiple cerebral infarctions | 120
brain MRI multiple cerebral infarctions | 120
POD 11 weaned to CPAP | 264
extubated | 264
POD 15 vital signs unstable | 360
catecholamines administration started | 360
panperitonitis confirmed | 360
gram (+) cocci on peritoneal culture | 360
POD 31 expired | 744
cardiac arrest | 744
septic shock | 744
