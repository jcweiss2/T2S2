39 years old | 0 | 0 
female | 0 | 0 
height 155 cm | 0 | 0 
weight 44.5 kg | 0 | 0 
mild dyspnea | 0 | 0 
adenoid cystic carcinoma in the carina | 0 | 0 
carinal resection | 0 | 360 
reconstruction | 0 | 360 
chest computed tomography | -24 | -24 
bronchoscopy | -24 | -24 
left mainstem bronchus obstruction | -24 | 0 
carina obstruction | -24 | 0 
right mainstem bronchus obstruction | -24 | 0 
internal diameter of RMB 11 mm | -24 | -24 
length of RMB 12 mm | -24 | -24 
length of distal LMB 20 mm | -24 | -24 
moderate obstructive pattern of pulmonary function test | -24 | -24 
forced expiratory volume in one second 1.88 liter | -24 | -24 
forced vital capacity 2.81 liter | -24 | -24 
ratio of forced expiratory volume in one second to forced vital capacity 67% | -24 | -24 
general anesthesia | 0 | 360 
target-controlled infusion of propofol | 0 | 360 
target-controlled infusion of remifentanil | 0 | 360 
rocuronium | 0 | 360 
tracheal intubation | 0 | 360 
right-sided double-lumen tube | 0 | 20 
right lateral position | 0 | 360 
left bronchi and vasculature dissection | 0 | 20 
thoracoscopic surgery | 0 | 20 
right OLV | 0 | 20 
arterial oxygen tension 462 mmHg | 20 | 20 
inspired oxygen fraction 1.0 | 0 | 360 
left thoracoscopic surgery | 20 | 40 
single-lumen endotracheal tube | 20 | 360 
bronchial blocker | 20 | 360 
left lateral position | 40 | 360 
right thoracotomy | 40 | 360 
peak airway pressure 28 cmH2O | 40 | 40 
tidal volume 300 ml | 40 | 40 
arterial oxygen tension 110 mmHg | 60 | 60 
left OLV | 40 | 360 
carinal resection | 60 | 360 
resection of LMB | 60 | 360 
insertion of sterile endotracheal tube into LMB | 60 | 360 
airway pressure 35 cmH2O | 60 | 60 
oxygen saturation by pulse oximetry 70% | 60 | 60 
resection of RMB | 60 | 360 
insertion of additional sterile endotracheal tube into RMB | 60 | 360 
differential bilateral lung ventilation | 60 | 360 
oxygen saturation by pulse oximetry 100% | 62 | 360 
removal of carina | 62 | 360 
anastomosis of RMB and trachea | 62 | 360 
no air leak in anastomotic site | 62 | 360 
removal of left endobronchial tube | 120 | 360 
non-dependent right OLV | 120 | 360 
low tidal volume 200-250 ml | 120 | 360 
airway pressure lower than 20 cmH2O | 120 | 360 
oxygen saturation by pulse oximetry below 80% | 120 | 120 
reinsertion of left endobronchial tube | 120 | 360 
two-lung ventilation | 120 | 360 
inspired oxygen fraction 1.0 | 120 | 360 
oxygen saturation by pulse oximetry 100% | 125 | 360 
right OLV | 125 | 360 
oxygen saturation by pulse oximetry below 90% | 128 | 128 
clamping of left pulmonary artery | 128 | 360 
ligation of left pulmonary artery | 128 | 360 
oxygen saturation by pulse oximetry 100% | 133 | 360 
removal of left endobronchial tube | 133 | 360 
closure of right thoracotomy | 133 | 360 
left thoracotomy | 180 | 360 
resection of left pulmonary artery and veins | 180 | 360 
left pneumonectomy | 180 | 360 
supine position | 360 | 360 
tracheal extubation | 360 | 360 
transfer to intensive care unit | 360 | 360 
discharge on 13th postoperative day | 780 | 780 
no complications | 780 | 780