23 years old | 0
male | 0
previous deceased-donor renal transplant | -43800
end-stage renal disease (ESRD) | -43800
membranoproliferative glomerulonephritis (MPGN) | -43800
tacrolimus | -43800
prednisone | -43800
constitutional symptoms | -336
intermittent fever | -336
fatigue | -336
blood pressure of 112/67 mmHg | 0
heart rate of 103 beats per minute | 0
pulse oximetry of 98% | 0
temperature of 37.1°C | 0
body mass index of 22.6 kg/m² | 0
S3 | 0
new-onset 3/6 holosystolic murmur | 0
scattered crackles | 0
mild peripheral edema | 0
COVID-19 PCR negative | 0
12-lead electrocardiogram with sinus tachycardia | 0
portable chest radiograph with pulmonary edema | 0
leukocytosis | 0
thrombocytosis | 0
normal hemoglobin | 0
mild acute kidney injury | 0
normal hepatic function panel | 0
normal coagulation studies | 0
elevated cardiac troponin | 0
elevated NT-proBNP | 0
elevated D-dimer | 0
hospitalized | 0
suspected infective endocarditis | 0
acute heart failure | 0
shifted to intensive care unit | 0
meropenem | 0
linezolid |-
levofloxacin | 0
fluconazole | 0
low-dose nitroglycerin | 0
furosemide infusions | 0
transthoracic echocardiogram with vegetation on mitral valve | 0
mitral valve perforation | 0
ruptured chordae tendinae | 0
torrential mitral regurgitation | 0
vegetation on aortic valve | 0
torrential aortic regurgitation | 0
repeat transthoracic echocardiogram with enlargement of vegetations | 72
deteriorating valve function | 72
positive Bartonella henselae IgM | 72
positive Coxiella burnetii IgM | 72
intravenous doxycycline | 72
intravenous gentamicin | 72
transesophageal echocardiogram with bicuspid aortic valve | 72
dual valve replacement | 168
aspirin | 168
warfarin | 168
uneventful postoperative course | 168
outpatient clinic follow-up at 10 days | 240
outpatient clinic follow-up at 1 month | 720
evaluated at 3 months post-discharge | 2160
no prosthetic valve endocarditis | 2160
no valve dysfunction | 2160
hydroxychloroquine therapy | 2160
clinically well | 2160
