40 years old | 0
    woman | 0
    presented to an outside emergency department (ED) | -48
    facial swelling | -48
    neck swelling | -48
    abdominal discomfort | -48
    tooth abscess | -72
    clindamycin | -72
    swelling of face worsened | 0
    swelling of neck worsened | 0
    endotracheal intubation | 0
    mechanical ventilation | 0
    CT scan neck | 0
    necrotizing fasciitis | 0
    soft tissue edema | 0
    gas formation | 0
    retropharyngeal abscess | 0
    tachycardic | 0
    tachypneic | 0
    blood pressure 89/41 mmHg | 0
    MAP 69 mmHg | 0
    WBC count 6.7 | 0
    H&H 12.5/37.2 | 0
    creatinine 1.8 | 0
    lactic acid 2.9 | 0
    central venous line placement | 0
    IV fluids 3 liters | 0
    transferred to ICU | 0
    necrotizing fasciitis | 0
    soft tissue abscess | 0
    progressing mediastinitis | 0
    fluid resuscitation | 0
    sedation on Versed | 0
    marked swelling of neck | 0
    rhonchorous breath sounds | 0
    severe sepsis | 0
    multiple organ dysfunction syndrome | 0
    deep soft tissue infection | 0
    intravenous Fentanyl | 0
    Sodium Chloride 1 liter | 0
    clindamycin | 0
    piperacillin-tazobactam | 0
    vancomycin | 0
    heparin | 0
    pantoprazole | 0
    Levophed infusion | 0
    ENT surgical debridement | 0
    packed submandibular incisions | 0
    packed anterior neck incisions | 0
    removed two teeth | 0
    right radial arterial line | 0
    CT chest | 24
    small pericardial effusion | 24
    moderate bilateral pleural effusions | 24
    loculation on left side | 24
    ground glass opacities | 24
    nodular consolidation | 24
    acute lung injury/ARDS | 24
    bilateral chest tubes | 24
    tracheostomy | 96
    PEG tube | 96
    pericardiocentesis | 240
    PICC line | 264
    culture neck wound | 264
    Clostridium subterminale | 264
    culture pleural fluid | 336
    Clostridium subterminale | 336
    sensitivity ampicillin-sulbactam | 336
    sensitivity cefoxitin | 336
    sensitivity meropenem | 336
    sensitivity metronidazole | 336
    sensitivity penicillin | 336
    full course piperacillin-tazobactam | 336
    maintenance enteral antibiotic therapy | 336
    chest tubes removed | 624
    discharged | 888
