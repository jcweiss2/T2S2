72 years old | 0
female | 0
admitted to the hospital | 0
bulging mass on her low abdomen | 0
ventral hernia repair | -120
severe abdominal pain | -120
septic shock | -120
exploratory laparotomy | -120
intestinal adhesions | -120
intraperitoneal contamination | -120
open drain system | -120
critical care | -120
systemic infection | -120
two EAFs | -96
well-controlled hypertension | 0
well-controlled diabetes | 0
no medical comorbidities | 0
no personal and family history | 0
physical examination | 0
bulging mass on her low abdomen | 0
no symptoms or signs of the intestinal obstruction | 0
laboratory examinations | 0
no abnormalities | 0
complete blood cell count | 0
cardiac markers | 0
coagulation profile | 0
abdominal computed tomography scan | 0
EAF on the midline of the abdomen | 0
fasting | 0
full caloric parenteral nutrition | 0
electrolyte repletion | 0
antacids | 0
octreotide | 0
frequent surgical wound dressing | 0
protection of the surrounding tissue from the enteric effluent | 0
vacuum-assisted closure dressings | 0
daily output of the EAFs consistently exceeded 1000 mL | 0
surrounding tissues severely contaminated by enteric effluent | 0
initiation of enteral nutrition | 0
output increased dramatically | 0
rubber drains inserted into the intestinal lumens | 24
fistula output decreased to < 500 mL/d | 24
endoscopic stent insertion | 48
expulsion of the inserted stents | 48
vascular grafts implanted | 768
enteric continuity restored | 768
anastomoses between the intestinal openings of each EAF and the vascular grafts | 768
no fistula output observed | 768
elemental EN began | 773
anastomoses not completely healed | 773
leakage after the initiation of elemental enteral feeding | 773
output remained < 300 mL/d | 773
patient became comfortable clinically and emotionally | 773
discharged from the hospital | 1056
VAC dressing management regularly at the outpatient department | 1056
EAF resection | 1344
involved intestines were the distal jejunum and sigmoid colon | 1344