48 years old| 0  
    male | 0  
    obese | 0  
    non-alcoholic steatohepatitis | 0  
    SARS-CoV-2 infection | 0  
    ground-glass pattern on thoracic CT | 0  
    positive nasopharyngeal swab test | 0  
    isolated in the Department of Infectious Diseases | 0  
    oseltamivir | 0  
    hydroxychloroquine | 0  
    broad-spectrum antibiotics | 0  
    endotracheal intubation | 72  
    invasive mechanical ventilation | 72  
    respiratory failure | 72  
    favipiravir | 72  
    rehabilitation program could not be implemented | 72  
    ARDS | 72  
    cardiopulmonary stability | 0  
    SARS-CoV-2 negativity confirmed | 0  
    in-bed positioning every 2 hours | 0  
    passive range of motion | 0  
    prone position 12-16 hours per day | 0  
    cytokine storm syndrome | 168  
    candidemia | 168  
    intravenous tocilizumab | 168  
    immune plasma | 168  
    intravenous high-dose glucocorticoids | 168  
    antifungal therapy | 168  
    clinical stability | 0  
    weaning | 0  
    controlled breathing techniques | 0  
    bronchial hygiene-airway clearance techniques | 0  
    home-based respiratory muscle exercise program | 0  
    threshold inspiratory muscle trainer device | 0  
    admitted to the inpatient clinic of PMR | 1704  
    weakness predominantly distal muscles of upper and lower extremities | 1704  
    right wrist drop | 1704  
    bilateral foot drop | 1704  
    symmetrical mild distal muscle atrophy | 1704  
    contractures of left hip | 1704  
    contractures of left knee | 1704  
    sacral decubitus ulcer | 1704  
    sensorimotor axonal peripheral neuropathy | 1704  
    cardiopulmonary functions could not be assessed | 1704  
    no respiratory function tests performed | 1704  
    thoracic CT no new findings | 1704  
    echocardiography no new findings | 1704  
    mild hypoalbuminemia | 1704  
    isolated low creatinine levels | 1704  
    ICU-AW originating from CIP | 1704  
    Mini-Mental State Examination score 25 | 1704  
    General Health Perception score 5 | 1704  
    Mental Health Perception score 0 | 1704  
    Physical Function score 0 | 1704  
    Functional Ambulation Category level 0 | 1704  
    MRC muscle strength score 30 | 1704  
    postural hypotensive attacks | 1704  
    tilt table training | 1704  
    active-assisted ROM | 1704  
    active ROM | 1704  
    isometric strength exercises | 1704  
    isotonic strength exercises | 1704  
    mobilization efforts | 1704  
    physical rehabilitation program 2 hours daily | 1704  
    physiotherapist accompaniment | 1704  
    methenolone enanthate 400 mg/week | 1704  
    neuromuscular electrical stimulation | 1704  
    collagen-containing dressing for sacral ulcer | 1704  
    walk with ankle-foot orthosis | 1704  
    walk with walker | 1704  
    improvement in MMSE score | 1704  
    improvement in SF-36 scores | 1704  
    hand grip strength measurements | 1704  
    pinch strength measurements | 1704  
    manual muscle testing using MRC scale | 1704  
    hand-held dynamometry | 1704  
    written informed consent obtained | 1704  
    early rehabilitation interventions | 1704  
    multidisciplinary team work | 1704  
    patient-specific rehabilitation plan | 1704  
    gradual progression of rehabilitation | 1704  
    passive ROM in admission period | 1704  
    passive cycling | 1704  
    electrical muscle stimulation | 1704  
    strengthening exercises | 1704  
    endurance exercises | 1704  
    balance exercises | 1704  
    occupational activities | 1704  
    methenolone enanthate use | 1704  
    tele-rehabilitation services discussed | 1704  
    home-based exercise programs explained | 1704  
    nutrition education for muscle remodeling | 1704  
    diet education for obesity prevention | 1704  
    hospital discharge | 1704  
    improved functional capacity | 1704  
    limited disability | 1704  
    no cardiopulmonary complications during rehabilitation | 1704  
    no exercise-induced desaturation | 1704  
    no spread risk of SARS-CoV-2 | 1704  
    no new cardiopulmonary findings | 1704  
    no heart failure | 1704  
    no heart valve pathologies | 1704  
    normal acute phase reactants | 1704  
    normal serum electrolytes | 1704  
    normal liver function tests | 1704  
    normal kidney function tests | 1704  
    secondary causes ruled out | 1704  
    favorable prognosis | 1704  
    improved quality of life | 1704  
    safe rehabilitation procedures | 1704  
    no increased mortality | 1704  
    no long-term complications | 1704  
    no neurological complications | 1704  
    no immune-mediated effects on myofibrils | 1704  
    no hyperglycemia | 1704  
    minimal sedation | 1704  
    no neuromuscular blockers | 1704  
    no barotrauma | 1704  
    no prolonged ICU stay | 1704  
    no subsequent development of obesity | 1704  
    no impaired lung function | 1704  
    no physiological impairment | 1704  
    no cognitive impairment | 1704  
    no mental impairment | 1704  
    no conflicts of interest | 1704  
    no financial support | 1704  
    discharged | 1704  

    