44 years old | 0
man | 0
transferred to our hospital | 0
intubated for hypoxia | -48
COVID-19-related pneumonia | -48
dry cough | -120
fever | -120
denied gastrointestinal symptoms | 0
denied myalgias | 0
denied dyspnea | 0
hypertension | 0
type II diabetes mellitus | 0
previous stroke secondary to left atrial thrombus | 0
outpatient treatment for diabetes | 0
metformin | 0
alogliptin | 0
serum glucose 222 mg/dL | 0
hemoglobin A1C not tested | 0
chest radiograph revealed patchy ground-glass opacities | 0
severe acute respiratory syndrome coronavirus 2 RT-PCR test positive | 0
human immunodeficiency virus antibody test negative | 0
white blood cell count 16.9 | 0
azithromycin | -48
ceftriaxone | -48
hydroxychloroquine | -48
developed worsening hypoxemia | -24
intubated | -24
received cefepime | -24
received vancomycin | -24
transferred to medical intensive care unit | 0
temperature 102.8°F | 0
blood pressure 138/77 mm Hg | 0
pulse 114 beats per minute | 0
respirations 16 | 0
oxygen saturation 95% | 0
mechanically ventilated | 0
weight 91 kilograms | 0
WBC 17.1 | 0
lactate dehydrogenase 570 | 0
C-reactive protein 328 | 0
ferritin 2043 | 0
d-dimer 0.74 | 0
interleukin-6 21 | 0
procalcitonin 5.59 | 0
vancomycin continued | 0
cefepime continued | 0
dexamethasone 20 mg/day | 72
methylprednisolone 40 mg | 168
cumulative dose equivalent to 717 mg prednisone | 168
QuantiFERON-TB Gold Plus test obtained | 96
QFT-Plus negative | 96
repeat specimen insufficient | 96
TCZ 400 mg intravenously | 96
afebrile | 120
WBC 24.9 | 168
temperature rose to 102°F | 192
piperacillin/tazobactam | 192
vancomycin | 192
self-extubation | 192
reintubation | 192
tracheal aspirate negative | 192
blood cultures negative | 192
clinical status improved | 192
fever resolution | 192
extubated | 384
BiPAP | 384
nasal cannula | 384
transferred to general medicine floor | 384
leukocytosis persisted | 384
temperature rose to 101.1°F | 528
WBC 14.7 | 528
left shift | 528
altered mental status | 528
treated with TZP | 528
fever persisted | 528
leukocytosis persisted | 528
vancomycin added | 576
blood cultures negative | 576
urine cultures negative | 576
fungal cultures negative | 576
serum galactomannan negative | 576
beta-d-glucan negative | 576
urinalysis negative | 576
chest radiograph revealed patchy infiltrates | 576
sputum Gram stain moderate Gram-positive cocci | 576
culture moderate growth Klebsiella pneumoniae | 576
TZP discontinued | 576
cefepime added | 576
fever persisted | 576
leukocytosis persisted | 576
sputum cultures negative | 576
CT scan chest and abdomen | 696
chest radiograph 1 day before CT scan | 672
meropenem | 696
caspofungin | 696
vancomycin | 696
metronidazole | 696
caspofungin discontinued | 768
voriconazole added | 768
leukocytosis | 768
intermittent fever | 768
sputum cultures negative | 768
CT scan chest | 840
blood cultures negative | 840
urine Legionella antigen negative | 840
serum galactomannan negative | 840
beta-d-glucan negative | 840
urine Histoplasma antigen negative | 840
Coccidioides IgG antibody negative | 840
repeat COVID-19 RT-PCR negative | 840
sputum smears positive for acid-fast bacilli | 840
MTB complex identified | 840
no rifampin resistance detected | 840
positive PPD test | 840
prior 3 months TB treatment | 840
born in Haiti | 840
travels to Haiti regularly | 840
antibiotics discontinued | 840
antifungal agents discontinued | 840
treated with isoniazid | 840
rifampin | 840
ethambutol | 840
pyrazinamide | 840
vitamin B6 | 840
oxygen saturation improved | 840
fever resolved | 840
leukocytosis resolved | 840
discharged | 864
serum glucose ranged 50-450 mg/dL | 864
45% serum glucose >180 | 864
pulmonary cavitary TB | 864
