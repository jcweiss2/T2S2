baby boy | 0
born by emergency cesarean section | 0
severe preeclampsia in the mother | -672
gestational week 25 6/7 | 0
birthweight 665 g | 0
intubated in the delivery room | 0
transferred to the neonatal intensive care unit | 0
mechanical ventilation | 0
total parenteral nutrition | 24
minimal enteral nutrition with breast milk | 24
delayed meconium passage | 48
abdominal distension | 48
increased gastric residuals | 48
necrotizing enterocolitis | 48
gastric free drainage | 144
broad-spectrum antibiotic therapy | 144
perforated NEC | 144
surgery | 144
short bowel syndrome | 168
thyroid screening tests | 336
low circulating free and total throxine | 336
low TSH | 336
high cortisol | 336
high serum total bilirubin level | 336
high direct reacting bilirubin | 336
enteral levothyroxine 5 µg/kg/day | 336
no response to treatment | 504
enteral levothyroxine 10 µg/kg/day | 504
poor absorption of the drug | 504
rectal levothyroxine 10 µg/kg/day | 576
increased fT4 levels | 624
decreased bilirubin levels | 624
died on postnatal 77th day | 1848
severe bronchopulmonary dysplasia | 1848
surgical NEC | 1848
short bowel syndrome | 1848
sepsis | 1848