38 years old | 0
female | 0
G4P3A0 L0 | 0
admitted to hospital | 0
unexplained fetal loss | -672
unexplained fetal loss | -1344
unexplained fetal loss | -2016
hypocellular bone marrow | -672
severe thrombocytopenia | -672
pregnancy induced hypertension (PIH) | -672
referred to Tertiary Care Center | -672
hemodynamically stable | 0
blood pressure 140/90 mmHg | 0
Tab. methyldopa 250 mg | -672
total leukocyte count 7200/μL | 0
hemoglobin (Hb) 8.5 g/dl | 0
hematocrit 22.6% | 0
platelet count 6000/mm3 | 0
blood group O negative | 0
pancytopenia | 0
bone marrow biopsy | 0
hypoplastic marrow | 0
Intrauterine growth retardation (IUGR) | 0
fetal well-being | 0
received 20 units of platelets | 0
received 2 units of whole blood | 0
oral prednisolone 10 mg tid | 0
oral hematinic | 0
antiplatelet antibody negative | 0
ANA negative | 0
antigen test for paroxysmal nocturnal hemoglobinopathies negative | 0
factor V mutation negative | 0
direct comb's test negative | 0
Fanconi anemia negative | 0
Hb electrophoresis normal | 0
leaking per vaginal | 24
Ultra sonography (USG) Doppler showed IUGR | 24
intermittent absent end diastolic flow | 24
posted for emergency lower segment cesarean section (LSCS) | 24
adequate units of blood arranged | 24
single donor platelets arranged | 24
fasting status confirmed | 24
high-risk written informed consent taken | 24
general anesthesia | 24
Electrocardiogram | 24
Oxygen saturation | 24
Non-invasive Blood Pressure monitors | 24
IV Nitroglycerine 60 μg | 24
IV metoprolol 1.5 mg | 24
6 units of platelets transfused | 24
IV Ranitidine 50 mg | 24
IV ondonsetron 4 mg | 24
IV glycopyrrolate 0.2 mg | 24
IV hydrocortisone 100 mg | 24
pre-oxygenated with 100% oxygen | 24
thiopentone sodium 300 mg | 24
tracheal intubation | 24
succinylcholine 100 mg | 24
IV xylocard 50 mg | 24
nitrous oxide-oxygen-vecuronium | 24
female infant weighing 960 g delivered | 24
poor Apgar scores | 24
shifted to neonatal intensive care unit (NICU) | 24
midazolam 1 mg | 24
fentanyl 100 μg | 24
stable hemodynamics intra-operatively | 24
total blood loss 1200 ml | 24
2 units of blood transfused | 24
10 units of platelets transfused | 24
neuromuscular blockade reversed | 24
trachea extubated | 24
shifted to Post-operative Anesthesia Care Unit (PACU) | 24
2 units of blood | 24
3 units of cryoprecipitates | 24
12 units of platelets | 24
prophylactic antibiotics | 24
IV cefuroxime 1.2 gm | 24
IV metronidazole 500 mg | 24
post-operative analgesia | 24
IV paracetamol 15 mg/kg | 24
post-operative persistent hypertension | 24
Nitroglycerine @ 0.5-1 μg/kg/h | 24
Labetalol 100 mg | 48
oral prednisolone 10 mg | 48
Hb 9.8 gm | 48
platelet count 28000/mm3 | 48
shifted to ward | 72
discharged from hospital | 240
followed-up in obstetric and hematology clinic | 240
planned for bone marrow transplant | 240