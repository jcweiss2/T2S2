18 years old | 0
male | 0
stabbed herself in the abdomen | 0
suicidal intent | 0
admitted to the emergency department | 0
blood pressure could not be measured | 0
pulseless electrical activity | 0
body temperature 35.0°C | 0
oxygen saturation 99% | 0
Glasgow Coma Scale score 3 | 0
agonal respiration | 0
wound on upper abdomen | 0
intra-abdominal fluid collection | 0
emergency thoracotomy | 0
aortic cross-clamping | 0
open cardiac massage | 0
epinephrine administered | 0
return of circulation | 0
hemodynamically unstable | 0
laparotomy | 0
injuries to the common hepatic and splenic arteries | 0
pancreas injury | 0
spleen injury | 0
liver injury | 0
ligation of the injured arteries | 0
distal pancreatectomy | 0
splenectomy | 0
liver sutured | 0
norepinephrine administered | 0
second-look surgery | 24
no signs of active bleeding | 24
no ischemic change | 24
no vasopressor requirement | 72
abdominal wall closure | 72
CT scan | 96
disruption of the celiac artery | 96
gastroduodenal artery arising from superior mesenteric artery | 96
gastroscopy | 120
patchy mucosal necrosis on the gastric upper body | 120
fever | 552
pain in the stomach | 552
white blood cell count 34,000/mm3 | 552
C reactive protein 13.4 mg/dL | 552
CT scan | 552
air in the gastric wall | 552
intra-abdominal free air | 552
emergency surgery | 552
necrosis of the stomach | 552
total gastrectomy with Roux-en-Y reconstruction | 552
histological findings of the stomach | 552
diffuse necrotic changes | 552
inflammatory cell infiltrations | 552
sepsis due to multidrug-resistant Pseudomonas aeruginosa infection | 696
disseminated intravascular coagulation | 696
death | 696