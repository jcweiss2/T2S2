65 years old | 0
male | 0
allergic rhinitis | 0
eczema | 0
dyslipidemia | 0
benign prostatic hyperplasia | 0
left eye blurring of vision | -26280
left visual field quadrantanopia | 0
no papilloedema | 0
no other neurological deficit | 0
pituitary macroadenoma | 0
low cortisol | 0
low growth hormone | 0
low testosterone | 0
TSH and excision of the tumor | 0
polyuria | 24
cranial diabetes insipidus | 24
desmopressin | 24
febrile | 168
tachypneic | 168
tachycardic | 168
minimal cough | 168
no neurological symptoms | 168
no cerebrospinal fluid rhinorrhea | 168
equal air entry in lungs | 168
no adventitious sound | 168
minimal perihilar haziness on chest X-ray | 168
WBC count 9000 cells/cm3 | 168
CRP 200 mg/L | 168
IV Tazosin started | 168
headache | 168
neck pain | 168
indecisive about lumbar puncture | 168
Glasgow Coma Scale drop (E4V5M6 to E3V3M5) | 216
pupils reactive 3/3 | 216
neck stiffness | 216
positive Kernig’s sign | 216
positive Brudzenski’s sign | 216
increased WBC to 14,000 cells/cm3 | 216
CRP >200 mg/L | 216
blood culture positive for E. meningoseptica | 216
septic shock | 216
intubated | 216
transferred to neurocritical care unit | 216
IV Meropenem started | 216
IV Ciprofloxacin started | 216
lumbar puncture | 216
CSF clear and yellowish | 216
CSF WBC increased 10 cells/mm3 | 216
CSF glucose 2.2 mmol/L | 216
CSF protein 0.57 g/L | 216
CSF culture positive for E. meningoseptica | 216
bacteremia diagnosis | 216
meningitis diagnosis | 216
no neurological improvement post antibiotics | 312
septic parameters improved | 312
contrast-enhanced CT brain | 312
superior sagittal sinus thrombosis | 312
SC clexane started | 312
tracheal aspirate culture grew Acinetobacter baumannii XDR | 312
IV Polymyxin B added | 312
IV Polymyxin completed for 14 days | 336
IV Meropenem completed for 14 days | 336
IV Ciprofloxacin completed for 14 days | 336
T. Levofloxacin started | 336
extubated | 408
culture and sensitivity completed | 336
venous sinus thrombosis resolving | 336
WBC 7000 cells/cm3 | 336
CRP negative | 336
full neurological recovery | 336
hospital discharge | 408
