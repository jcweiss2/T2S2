86 years old | 0
overweight | 0
female | 0
appendectomy | -51600
implantation of heart pacemaker | -8760
severe abdominal pain | -24
nausea | -24
vomiting | -24
dehydration | 0
tenderness | 0
elevation of pancreatic enzymes | 0
elevated serum amylase | 0
elevated urinary amylase | 0
elevated serum lipase | 0
elevated glucose level | 0
normal serum C-reactive protein level | 0
normal serum white blood cell count | 0
marginal dilatation of the common bile duct | 0
thin-walled gallbladder | 0
excessive bowel gas | 0
admitted to the surgery department | 0
strict diet | 0
intravenous hydration | 0
analgesic treatment | 0
persistent severe abdominal pain | 12
hypotension | 12
oliguria | 12
elevated serum C-reactive protein level | 12
decreased serum white blood cell count | 12
high percentage of neutrophils | 12
increased serum aspartate aminotransferase | 12
increased serum alanine aminotransferase | 12
computed tomography | 16
free gas in the peritoneal cavity | 16
free gas in the retroperitoneum | 16
perforated duodenal diverticulum | 16
emergency surgery | 16
perforation of the duodenum ruled out | 16
gangrenous gallbladder | 16
free fluid of purulent character | 16
cholecystectomy | 16
peritoneal cavity lavage | 16
drainage | 16
gas in the gallbladder wall | 16
gas in the pancreatic parenchyma | 16
pneumobilia | 16
penetration of gas into abdominal wall | 16
emphysematous cholecystitis | 16
gangrenous pancreatitis | 16
retroperitoneal gangrene | 16
septic shock | 24
multiorgan failure | 24
increased procalcitonin | 24
increased C-reactive protein | 24
increased D-dimer | 24
increased lactate dehydrogenase | 24
increased creatine phosphokinase | 24
increased myoglobin | 24
increased troponin | 24
decreased red blood cell count | 24
decreased haemoglobin level | 24
relaparotomy | 24
cardiac arrest | 24
death | 24