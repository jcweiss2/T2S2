61 years old | 0
female | 0
white | 0
Ashkenazi Jewish descent | 0
admitted to the hospital | 0
nausea | -192
vomiting | -192
fever | -192
edema | -192
splenomegaly | -192
palpable axillary lymph nodes | -192
mild anemia | 0
thrombocytopenia | 0
hypoalbuminemia | 0
elevated CRP | 0
elevated alkaline phosphatase | 0
elevated GGT | 0
elevated IL-6 | 0
lymphoid hyperplasia | 0
lymph node biopsy | 0
bone marrow biopsy | 0
renal biopsy | 0
PET-CT scan | 0
bilateral pleural effusion | 0
retroperitoneal lymph node enlargement | 0
admitted to ICU | 168
worsening of anasarca | 168
worsening of renal function | 168
multiple organ failure | 168
mechanical ventilation | 168
CRRT | 168
diagnosis of TAFRO syndrome | 432
methylprednisolone started | 432
tocilizumab started | 432
rituximab started | 432
improvement in respiratory status | 600
improvement in hemodynamic status | 600
intermittent hemodialysis | 936
discharged from ICU | 1104
discharged from hospital | 2160
TAFRO syndrome | 0
anasarca | 0
organomegaly | 0
bone marrow fibrosis | 0
renal failure | 0
thrombocytopenia | 0
fever | -192
renal thrombotic microangiopathy | 0
mesangial expansion | 0
duplication of capillary basal membrane | 0
elevated IL-6 | 0
tocilizumab | 432
rituximab | 432
methylprednisolone | 432
steroids | 432
anti-IL-6 antibodies | 432
complete resolution of anasarca | 2160
complete resolution of organomegaly | 2160
normalization of hemoglobin | 2160
normalization of platelet count | 2160
decrease in IL-6 levels | 2160