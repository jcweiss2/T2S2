66 years old | 0
male | 0
SARS-CoV-2 infection | -1464
septic shock | -1464
hemodynamic instability | -1464
orotracheal intubation | -1464
pulmonary insufficiency | -1464
renal failure | -1464
admitted to the hospital | 0
arterial hypertension | 0
moderate alcoholism | 0
coronary disease | 0
Dieulafoy gastric lesion | 0
esophageal ulcers | 0
cytomegalovirus infection | 0
hepatomegaly | 0
blood transfusions | 0
antibiotics | 0
corticosteroids | 0
ganciclovir | 0
acute kidney injury | 0
hemodialysis | 0
hemodynamic improvement | 0
pulmonary improvement | 0
renal improvement | 0
CMV treatment | 0
cholestatic enzymes increase | 0
metabolic markers negative | 0
genetic markers negative | 0
autoimmune hepatic disease antibodies negative | 0
serologies negative | 0
PCRs for viruses negative | 0
immunoglobulin levels normal | 0
MRCP findings | 0
biliary cast | 0
serum ammonia >250 | 0
neurological symptoms | 0
sodium benzoate | 0
ursodeoxycholic acid | 0
serum ammonia decrease | 24
neurological function partial recovery | 24
liver function deterioration | 24
liver biopsy | 0
bile ductular reaction | 0
cholangiocyte injury | 0
inflammatory infiltrate | 0
biliary infarctions | 0
marked cholestasis | 0
portal fibrosis | 0
degenerative cholangiocyte injury | 0
cholangiocyte cytoplasmic vacuolization | 0
degenerative changes | 0
no thrombosis | 0
no bile duct dilatation | 0
no chronic liver disease | 0
no alcoholic hepatitis | 0
AST peak | 0
ALT peak | 0
bilirubin increase | 0
cholestatic liver enzymes increase | 0
hyperbilirubinemia | 0
no intrahepatic microangiopathy | 0
liver transplantation not performed | 24
discharged | 2928
