29 years old | 0
    female | 0
    pregnant | 0
    33-week 5-day period of gestation | 0
    fever | -144
    chills | -144
    nonproductive cough | -144
    breathlessness | -24
    continuous high-grade fever (103°F) | -144
    chills | -144
    rigor | -144
    no evening rise | -144
    no weight loss | -144
    dry nonproductive cough | -144
    running nose | -144
    sore throat | -144
    postnasal drip | -144
    sudden onset breathlessness | -24
    breathlessness progressed to symptomatic at rest | -24
    breathlessness aggravated with mild exertion | -24
    malaise | -144
    body ache | -144
    lethargy | -144
    weakness | -144
    tachycardia (108/min) | 0
    tachypnea (RR 26/min) | 0
    blood pressure 140/92 mmHg | 0
    SPO2 90%-92% at room air | 0
    SPO2 98% with oxygen supplementation | 0
    bilateral crackles | 0
    bilateral nonhomogeneous opacity on chest X-ray | 0
    admitted to respiratory ICU | 0
    suspicion of viral pneumonia | 0
    suspicion of ARDS | 0
    confirmed H1N1 infection | 0
    started oseltamivir 75 mg BD | 0
    started azithromycin 500 mg TDS | 0
    started paracetamol 15 mg/kg TDS | 0
    urgent consultation for termination of pregnancy at 34 weeks | 0
    steroid prophylaxis for fetal lung maturity | 0
    THRIVE therapy initiation | 0
    hemodynamic monitoring | 0
    high-risk consent for surgery | 0
    health-care professionals briefed | 0
    personal protection worn | 0
    wheeled to OT with Airvo™ 2 device | 0
    oxygen saturation 98% | 0
    RR 24/min | 0
    FiO2 0.5 | 0
    ABG pH 7.38 | 0
    ABG PCO2 38 mmHg | 0
    ABG PO2 110 mmHg | 0
    ABG HCO3 22 mmol/L | 0
    standard monitoring | 0
    spinal anesthesia administered | 0
    NIV (ResMed) standby | 0
    emergency intubation preparations | 0
    spinal anesthesia in sitting position | 0
    bupivacaine heavy 0.5% given | 0
    supine with left tilt | 0
    head raised with pillows | 0
    high-flow oxygen continued | 0
    block level confirmed to T4 | 0
    surgery started | 0
    two healthy female infants born | 0
    uterotonics titrated | 0
    continuous intraoperative monitoring | 0
    IV plasmalyte 500 ml administered | 0
    RR 24-26/min during surgery | 0
    bilateral transversus abdominis plane block | 0
    postoperative breathlessness | 24
    RR increased to 40/min | 24
    SpO2 90% | 24
    placed on NIV | 24
    furosemide 40 mg IV | 24
    shifted to ICU | 24
    ABG pH 7.30 | 24
    ABG PCO2 48 mmHg | 24
    ABG PO2 68 mmHg | 24
    ABG HCO3 19 mmol/L | 24
    RR reduced to 22/min | 48
    ABG pH 7.36 | 48
    ABG PCO2 38 mmHg | 48
    ABG PO2 98 mmHg | 48
    ABG HCO3 20 mmol/L | 48
    weaned off NIV | 48
    favorable outcome for mother | 48
    favorable outcome for child | 48

