56 years old | 0 | 0 
female | 0 | 0 
admitted to the hospital | 0 | 0 
history of weakness | -720 | 0 
numbness and weakness in lower extremities | -720 | -672 
numbness and weakness progressed to hands and neck | -672 | -624 
presumptive diagnosis of Guillain-Barré syndrome (GBS) | -720 | -624 
type 2 diabetes mellitus | 0 | 0 
hypertension | 0 | 0 
necrotizing pancreatitis due to gallstones | -8760 | -8760 
severe protein-calorie malnutrition | -8760 | -168 
total parenteral nutrition (TPN) | -8760 | -168 
discontinuation of TPN | -168 | -168 
return to normal diet | -168 | 0 
lumbar puncture | 0 | 0 
albuminocytologic dissociation in cerebrospinal fluid (CSF) | 0 | 0 
brain magnetic resonance imaging (MRI) scan | 0 | 0 
small vessel ischemic changes | 0 | 0 
intravenous immunoglobulin (IVIG) treatment | 0 | 120 
worsening pancytopenia | 120 | 120 
encephalopathy | 120 | 120 
transfer to specialist center | 120 | 120 
hypotensive | 120 | 120 
unresponsive to verbal stimuli | 120 | 120 
minimally responsive to painful stimuli | 120 | 120 
Glasgow Coma Scale (GCS) score of 6 | 120 | 120 
anasarcic | 120 | 120 
flaccid paralysis of all four extremities | 120 | 120 
malnourished and septic state | 120 | 120 
calcium of 6.7 mg/dL | 120 | 120 
hemoglobin of 9.4 g/dL | 120 | 120 
white cell count of 2.1×10^9/L | 120 | 120 
phosphorus of 1.1 mg/dL | 120 | 120 
creatinine <0.2 mg/dL | 120 | 120 
albumin <1.5 gm/dL | 120 | 120 
lactate of 4 mmol/L | 120 | 120 
nutritional risk screening (NRS-2002) score of 5 | 120 | 120 
malnutrition universal screening (MUST) score of 5 | 120 | 120 
intubation | 120 | 120 
resuscitation with intravenous fluids | 120 | 120 
intravenous infusion of norepinephrine | 120 | 168 
meropenem treatment | 120 | 168 
vancomycin treatment | 120 | 168 
anidulafungin treatment | 120 | 168 
empirical treatment with high-dose intravenous thiamine | 120 | 336 
electroencephalogram (EEG) | 168 | 168 
diffuse slow waves consistent with severe metabolic encephalopathy | 168 | 168 
brain MRI scan | 168 | 168 
hyperintensity of bilateral medial thalamus | 168 | 168 
serum thiamine level of 104 nmol/L | 168 | 168 
improvement in mental status | 192 | 192 
ability to understand simple commands | 192 | 192 
discontinuation of norepinephrine and antimicrobial treatment | 192 | 192 
resolution of hemodynamic stability | 192 | 192 
negative blood and urine cultures | 192 | 192 
extubation | 120 | 120 
electromyography (EMG) | 168 | 168 
severe sensorimotor polyneuropathy | 168 | 168 
improvement in mentation and weakness | 192 | 336 
transfer out of intensive care unit (ICU) | 336 | 336 
discharge | 336 | 336 
thiamine supplementation | 120 | 336 
dry beriberi | 120 | 336 
Wernicke’s encephalopathy | 168 | 336 
ascending neuropathy | -720 | 0 
paralysis | -720 | 0 
autonomic instability | 120 | 120 
cardiomyopathy | 0 | 0 
cardiomegaly | 0 | 0 
dyspnea | 0 | 0 
peripheral edema | 0 | 0 
shoshin beriberi | 0 | 0 
cardiogenic shock | 0 | 0 
lactic acidosis | 0 | 0 
multi-organ failure | 0 | 0 
altered mental status | 120 | 120 
ataxia | 120 | 120 
ocular symptoms | 120 | 120 
irreversible cognitive impairment | 0 | 0 
axonal abnormalities | 0 | 0 
impaired acetylcholine transmission | 0 | 0 
ataxia | 0 | 0 
areflexia | 0 | 0 
painful sensory or sensorimotor polyneuropathy | 0 | 0 
muscle weakness | 0 | 0 
Guillain-Barré syndrome (GBS) | -720 | 120 
acute inflammatory demyelinating polyradiculoneuropathy (AIDP) | -720 | 120 
infection | 0 | 0 
electromyography | 168 | 168 
nerve histology | 0 | 0 
axonal degeneration | 0 | 0 
demyelination | 0 | 0 
albuminocytologic dissociation | 0 | 0 
chronic inflammatory demyelinating polyneuropathy (CIDP) | 0 | 0 
critical illness myopathy | 120 | 120 
critical illness polyneuropathy | 120 | 120 
sepsis | 120 | 120 
encephalopathy | 120 | 120 
delirium | 120 | 120 
mechanical ventilation | 120 | 120 
neuromuscular disorders | 0 | 0 
primary neuromuscular disorders | 0 | 0 
thiamine deficiency | -720 | 336 
beriberi | -720 | 336 
malabsorption | 0 | 0 
alcohol abuse | 0 | 0 
anorexia nervosa | 0 | 0 
dieting | 0 | 0 
bariatric surgery | 0 | 0 
diarrhea | 0 | 0 
celiac disease | 0 | 0 
tropical sprue | 0 | 0 
dysentery | 0 | 0 
burns | 0 | 0 
pregnancy | 0 | 0 
dialysis | 0 | 0 
malignancy | 0 | 0 
thiamine supplementation | 120 | 336 
high-dose intravenous thiamine | 120 | 336 
magnetic resonance imaging (MRI) | 168 | 168 
electrophysiological studies | 168 | 168 
neuropathy | 0 | 0 
weakness | 0 | 0 
cardiomyopathy | 0 | 0 
autonomic instability | 120 | 120 
thiamine deficiency resulting beriberi | -720 | 336 
Guillain-Barré syndrome (GBS) | -720 | 120 
acute inflammatory demyelinating polyneuropathy (AIDP) | -720 | 120 
dry beriberi | 120 | 336 
Wernicke’s encephalopathy | 168 | 336 
thiamine levels | 168 | 168 
thiamine repletion | 120 | 336 
intravenous thiamine | 120 | 336 
thiamine therapy | 120 | 336 
thiamine deficiency-associated neuropathy | 0 | 0 
GBS treatment | -720 | 120 
IVIG therapy | 0 | 120 
thiamine supplementation | 120 | 336 
neurologic symptoms | 0 | 0 
neurologic function | 192 | 336 
encephalopathy | 120 | 120 
ascending lower extremity weakness | -720 | 0 
cerebrospinal fluid (CSF) findings | 0 | 0 
intravenous immunoglobulin (IVIG) treatment | 0 | 120 
thiamine supplementation | 120 | 336 
central neurologic function | 192 | 336 
peripheral neurologic function | 192 | 336 
recovery | 192 | 336 
thiamine deficiency | -720 | 336 
beriberi | -720 | 336 
Guillain-Barré syndrome (GBS) | -720 | 120 
mimic | 0 | 0 
case reports | 0 | 0 
thiamine levels | 168 | 168 
thiamine repletion | 120 | 336 
thiamine therapy | 120 | 336 
thiamine deficiency-associated neuropathy | 0 | 0 
GBS treatment | -720 | 120 
IVIG therapy | 0 | 120 
thiamine supplementation | 120 | 336 
neurologic symptoms | 0 | 0 
neurologic function | 192 | 336 
encephalopathy | 120 | 120 
ascending lower extremity weakness | -720 | 0 
cerebrospinal fluid (CSF) findings | 0 | 0 
intravenous immunoglobulin (IVIG) treatment | 0 | 120 
thiamine supplementation | 120 | 336 
central neurologic function | 192 | 336 
peripheral neurologic function | 192 | 336 
recovery | 192 | 336 
thiamine deficiency | -720 | 336 
beriberi | -720 | 336 
Guillain-Barré syndrome (GBS) | -720 | 120 
mimic | 0 | 0 
case reports | 0 | 0 
thiamine levels | 168 | 168 
thiamine repletion | 120 | 336 
thiamine therapy | 120 | 336 
thiamine deficiency-associated neuropathy | 0 | 0 
GBS treatment | -720 | 120 
IVIG therapy | 0 | 120 
thiamine supplementation | 120 | 336 
neurologic symptoms | 0 | 0 
neurologic function | 192 | 336 
encephalopathy | 120 | 120 
ascending lower extremity weakness | -720 | 0 
cerebrospinal fluid (CSF) findings | 0 | 0 
intravenous immunoglobulin (IVIG) treatment | 0 | 120 
thiamine supplementation | 120 | 336 
central neurologic function | 192 | 336 
peripheral neurologic function | 192 | 336 
recovery | 192 | 336 
thiamine deficiency | -720 | 336 
beriberi | -720 | 336 
Guillain-Barré syndrome (GBS) | -720 | 120 
mimic | 0 | 0 
case reports | 0 | 0 
thiamine levels | 168 | 168 
thiamine repletion | 120 | 336 
thiamine therapy | 120 | 336 
thiamine deficiency-associated neuropathy | 0 | 0 
GBS treatment | -720 | 120 
IVIG therapy | 0 | 120 
thiamine supplementation | 120 | 336 
neurologic symptoms | 0 | 0 
neurologic function | 192 | 336 
encephalopathy | 120 | 120 
ascending lower extremity weakness | -720 | 0 
cerebrospinal fluid (CSF) findings | 0 | 0 
intravenous immunoglobulin (IVIG) treatment | 0 | 120 
thiamine supplementation | 120 | 336 
central neurologic function | 192 | 336 
peripheral neurologic function | 192 | 336 
recovery | 192 | 336 
thiamine deficiency | -720 | 336 
beriberi | -720 | 336 
Guillain-Barré syndrome (GBS) | -720 | 120 
mimic | 0 | 0 
case reports | 0 | 0 
thiamine levels | 168 | 168 
thiamine repletion | 120 | 336 
thiamine therapy | 120 | 336 
thiamine deficiency-associated neuropathy | 0 | 0 
GBS treatment | -720 | 120 
IVIG therapy | 0 | 120 
thiamine supplementation | 120 | 336 
neurologic symptoms | 0 | 0 
neurologic function | 192 | 336 
encephalopathy | 120 | 120 
ascending lower extremity weakness | -720 | 0 
cerebrospinal fluid (CSF) findings | 0 | 0 
intravenous immunoglobulin (IVIG) treatment | 0 | 120 
thiamine supplementation | 120 | 336 
central neurologic function | 192 | 336 
peripheral neurologic function | 192 | 336 
recovery | 192 | 336 
thiamine deficiency | -720 | 336 
beriberi | -720 | 336 
Guillain-Barré syndrome (GBS) | -720 | 120 
mimic | 0 | 0 
case reports | 0 | 0 
thiamine levels | 168 | 168 
thiamine repletion | 120 | 336 
thiamine therapy | 120 | 336 
thiamine deficiency-associated neuropathy | 0 | 0 
GBS treatment | -720 | 120 
IVIG therapy | 0 | 120 
thiamine supplementation | 120 | 336 
neurologic symptoms | 0 | 0 
neurologic function | 192 | 336 
encephalopathy | 120 | 120 
ascending lower extremity weakness | -720 | 0 
cerebrospinal fluid (CSF) findings | 0 | 0 
intravenous immunoglobulin (IVIG) treatment | 0 | 120 
thiamine supplementation | 120 | 336 
central neurologic function | 192 | 336 
peripheral neurologic function | 192 | 336 
recovery | 192 | 336 
thiamine deficiency | -720 | 336 
beriberi | -720 | 336 
Guillain-Barré syndrome (GBS) | -720 | 120 
mimic | 0 | 0 
case reports | 0 | 0 
thiamine levels | 168 | 168 
thiamine repletion | 120 | 336 
thiamine therapy | 120 | 336 
thiamine deficiency-associated neuropathy | 0 | 0 
GBS treatment | -720 | 120 
IVIG therapy | 0 | 120 
thiamine supplementation | 120 | 336 
neurologic symptoms | 0 | 0 
neurologic function | 192 | 336 
encephalopathy | 120 | 120 
ascending lower extremity weakness | -720 | 0 
cerebrospinal fluid (CSF) findings | 0 | 0 
intravenous immunoglobulin (IVIG) treatment | 0 | 120 
thiamine supplementation | 120 | 336 
central neurologic function | 192 | 336 
peripheral neurologic function | 192 | 336 
recovery | 192 | 336 
thiamine deficiency | -720 | 336 
beriberi | -720 | 336 
Guillain-Barré syndrome (GBS) | -720 | 120 
mimic | 0 | 0 
case reports | 0 | 0 
thiamine levels | 168 | 168 
thiamine repletion | 120 | 336 
thiamine therapy | 120 | 336 
thiamine deficiency-associated neuropathy | 0 | 0 
GBS treatment | -720 | 120 
IVIG therapy | 0 | 120 
thiamine supplementation | 120 | 336 
neurologic symptoms | 0 | 0 
neurologic function | 192 | 336 
encephalopathy | 120 | 120 
ascending lower extremity weakness | -720 | 0 
cerebrospinal fluid (CSF) findings | 0 | 0 
intravenous immunoglobulin (IVIG) treatment | 0 | 120 
thiamine supplementation | 120 | 336 
central neurologic function | 192 | 336 
peripheral neurologic function | 192 | 336 
recovery | 192 | 336 
thiamine deficiency | -720 | 336 
beriberi | -720 | 336 
Guillain-Barré syndrome (GBS) | -720 | 120 
mimic | 0 | 0 
case reports | 0 | 0 
thiamine levels | 168 | 168 
thiamine repletion | 120 | 336 
thiamine therapy | 120 | 336 
thiamine deficiency-associated neuropathy | 0 | 0 
GBS treatment | -720 | 120 
IVIG therapy | 0 | 120 
thiamine supplementation | 120 | 336 
neurologic symptoms | 0 | 0 
neurologic function | 192 | 336 
encephalopathy | 120 | 120 
ascending lower extremity weakness | -720 | 0 
cerebrospinal fluid (CSF) findings | 0 | 0 
intravenous immunoglobulin (IVIG) treatment | 0 | 120 
thiamine supplementation | 120 | 336 
central neurologic function | 192 | 336 
peripheral neurologic function | 192 | 336 
recovery | 192 | 336 
thiamine deficiency | -720 | 336 
beriberi | -720 | 336 
Guillain-Barré syndrome (GBS) | -720 | 120 
mimic | 0 | 0 
case reports | 0 | 0 
thiamine levels | 168 | 168 
thiamine repletion | 120 | 336 
thiamine therapy | 120 | 336 
thiamine deficiency-associated neuropathy | 0 | 0 
GBS treatment | -720 | 120 
IVIG therapy | 0 | 120 
thiamine supplementation | 120 | 336 
neurologic symptoms | 0 | 0 
neurologic function | 192 | 336 
encephalopathy | 120 | 120 
ascending lower extremity weakness | -720 | 0 
cerebrospinal fluid (CSF) findings | 0 | 0 
intravenous immunoglobulin (IVIG) treatment | 0 | 120 
thiamine supplementation | 120 | 336 
central neurologic function | 192 | 336 
peripheral neurologic function | 192 | 336 
recovery | 192 | 336 
thiamine deficiency | -720 | 336 
beriberi | -720 | 336 
Guillain-Barré syndrome (GBS) | -720 | 120 
mimic | 0 | 0 
case reports | 0 | 0 
thiamine levels | 168 | 168 
thiamine repletion | 120 | 336 
thiamine therapy | 120 | 336 
thiamine deficiency-associated neuropathy | 0 | 0 
GBS treatment | -720 | 120 
IVIG therapy | 0 | 120 
thiamine supplementation | 120 | 336 
neurologic symptoms | 0 | 0 
neurologic function | 192 | 336 
encephalopathy | 120 | 120 
ascending lower extremity weakness | -720 | 0 
cerebrospinal fluid (CSF) findings | 0 | 0 
intravenous immunoglobulin (IVIG) treatment | 0 | 120 
thiamine supplementation | 120 | 336 
central neurologic function | 192 | 336 
peripheral neurologic function | 192 | 336 
recovery | 192 | 336 
thiamine deficiency | -720 | 336 
beriberi | -720 | 336 
Guillain-Barré syndrome (GBS) | -720 | 120 
mimic | 0 | 0 
case reports | 0 | 0 
thiamine levels | 168 | 168 
thiamine repletion | 120 | 336 
thiamine therapy | 120 | 336 
thiamine deficiency-associated neuropathy | 0 | 0 
GBS treatment | -720 | 120 
IVIG therapy | 0 | 120 
thiamine supplementation | 120 | 336 
neurologic symptoms | 0 | 0 
neurologic function | 192 | 336 
encephalopathy | 120 | 120 
ascending lower extremity weakness | -720 | 0 
cerebrospinal fluid (CSF) findings | 0 | 0 
intravenous immunoglobulin (IVIG) treatment | 0 | 120 
thiamine supplementation | 120 | 336 
central neurologic function | 192 | 336 
peripheral neurologic function | 192 | 336 
recovery | 192 | 336 
thiamine deficiency | -720 | 336 
beriberi | -720 | 336 
Guillain-Barré syndrome (GBS) | -720 | 120 
mimic | 0 | 0 
case reports | 0 | 0 
thiamine levels | 168 | 168 
thiamine repletion | 120 | 336 
thiamine therapy | 120 | 336 
thiamine deficiency-associated neuropathy | 0 | 0 
GBS treatment | -720 | 120 
IVIG therapy | 0 | 120 
thiamine supplementation | 120 | 336 
neurologic symptoms | 0 | 0 
neurologic function | 192 | 336 
encephalopathy | 120 | 120 
ascending lower extremity weakness | -720 | 0 
cerebrospinal fluid (CSF) findings | 0 | 0 
intravenous immunoglobulin (IVIG) treatment | 0 | 120 
thiamine supplementation | 120 | 336 
central neurologic function | 192 | 336 
peripheral neurologic function | 192 | 336 
recovery | 192 | 336 
thiamine deficiency | -720 | 336 
beriberi | -720 | 336 
Guillain-Barré syndrome (GBS) | -720 | 120 
mimic | 0 | 0 
case reports | 0 | 0 
thiamine levels | 168 | 168 
thiamine repletion | 120 | 336 
thiamine therapy | 120 | 336 
thiamine deficiency-associated neuropathy | 0 | 0 
GBS treatment | -720 | 120 
IVIG therapy | 0 | 120 
thiamine supplementation | 120 | 336 
neurologic symptoms | 0 | 0 
neurologic function | 192 | 336 
encephalopathy | 120 | 120 
ascending lower extremity weakness | -720 | 0 
cerebrospinal fluid (CSF) findings | 0 | 0 
intravenous immunoglobulin (IVIG) treatment | 0 | 120 
thiamine supplementation | 120 | 336 
central neurologic function | 192 | 336 
peripheral neurologic function | 192 | 336 
recovery | 192 | 336 
thiamine deficiency | -720 | 336 
beriberi | -720 | 336 
Guillain-Barré syndrome (GBS) | -720 | 120 
mimic | 0 | 0 
case reports | 0 | 0 
thiamine levels | 168 | 168 
thiamine repletion | 120 | 336 
thiamine therapy | 120 | 336 
thiamine deficiency-associated neuropathy | 0 | 0 
GBS treatment | -720 | 120 
IVIG therapy | 0 | 120 
thiamine supplementation | 120 | 336 
neurologic symptoms | 0 | 0 
neurologic function | 192 | 336 
encephalopathy | 120 | 120 
ascending lower extremity weakness | -720 | 0 
cerebrospinal fluid (CSF) findings | 0 | 0 
intravenous immunoglobulin (IVIG) treatment | 0 | 120 
thiamine supplementation | 120 | 336 
central neurologic function | 192 | 336 
peripheral neurologic function | 192 | 336 
recovery | 192 | 336 
thiamine deficiency | -720 | 336 
beriberi | -720 | 336 
Guillain-Barré syndrome (GBS) | -720 | 120 
mimic | 0 | 0 
case reports | 0 | 0 
thiamine levels | 168 | 168 
thiamine repletion | 120 | 336 
thiamine therapy | 120 | 336 
thiamine deficiency-associated neuropathy | 0 | 0 
GBS treatment | -720 | 120 
IVIG therapy | 0 | 120 
thiamine supplementation | 120 | 336 
neurologic symptoms | 0 | 0 
neurologic function | 192 | 336 
encephalopathy | 120 | 120 
ascending lower extremity weakness | -720 | 0 
cerebrospinal fluid (CSF) findings | 0 | 0 
intravenous immunoglobulin (IVIG) treatment | 0 | 120 
thiamine supplementation | 120 | 336 
central neurologic function | 192 | 336 
peripheral neurologic function | 192 | 336 
recovery | 192 | 336 
thiamine deficiency | -720 | 336 
beriberi | -720 | 336 
Guillain-Barré syndrome (GBS) | -720 | 120 
mimic | 0 | 0 
case reports | 0 | 0 
thiamine levels | 168 | 168 
thiamine repletion | 120 | 336 
thiamine therapy | 120 | 336 
thiamine deficiency-associated neuropathy | 0 | 0 
GBS treatment | -720 | 120 
IVIG therapy | 0 | 120 
thiamine supplementation | 120 | 336 
neurologic symptoms | 0 | 0 
neurologic function | 192 | 336 
encephalopathy | 120 | 120 
ascending lower extremity weakness | -720 | 0 
cerebrospinal fluid (CSF) findings | 0 | 0 
intravenous immunoglobulin (IVIG) treatment | 0 | 120 
thiamine supplementation | 120 | 336 
central neurologic function | 192 | 336 
peripheral neurologic function | 192 | 336 
recovery | 192 | 336 
thiamine deficiency | -720 | 336 
beriberi | -720 | 336 
Guillain-Barré syndrome (GBS) | -720 | 120 
mimic | 0 | 0 
case reports | 0 | 0 
thiamine levels | 168 | 168 
thiamine repletion | 120 | 336 
thiamine therapy | 120 | 336 
thiamine deficiency-associated neuropathy | 0 | 0 
GBS treatment | -720 | 120 
IVIG therapy | 0 | 120 
thiamine supplementation | 120 | 336 
neurologic symptoms | 0 | 0 
neurologic function | 192 | 336 
encephalopathy | 120 | 120 
ascending lower extremity weakness | -720 | 0 
cerebrospinal fluid (CSF) findings | 0 | 0 
intravenous immunoglobulin (IVIG) treatment | 0 | 120 
thiamine supplementation | 120 | 336 
central neurologic function | 192 | 336 
peripheral neurologic function | 192 | 336 
recovery | 192 | 336 
thiamine deficiency | -720 | 336 
beriberi | -720 | 336 
Guillain-Barré syndrome (GBS) | -720 | 120 
mimic | 0 | 0 
case reports | 0 | 0 
thiamine levels | 168 | 168 
thiamine repletion | 120 | 336 
thiamine therapy | 120 | 336 
thiamine deficiency-associated neuropathy | 0 | 0 
GBS treatment | -720 | 120 
IVIG therapy | 0 | 120 
thiamine supplementation | 120 | 336 
neurologic symptoms | 0 | 0 
neurologic function | 192 | 336 
encephalopathy | 120 | 120 
ascending lower extremity weakness | -720 | 0 
cerebrospinal fluid (CSF) findings | 0 | 0 
intravenous immunoglobulin (IVIG) treatment | 0 | 120 
thiamine supplementation | 120 | 336 
central neurologic function | 192 | 336 
peripheral neurologic function | 192 | 336 
recovery | 192 | 336 
thiamine deficiency | -720 | 336 
beriberi | -720 | 336 
Guillain-Barré syndrome (GBS) | -720 | 120 
mimic | 0 | 0 
case reports | 0 | 0 
thiamine levels | 168 | 168 
thiamine repletion | 120 | 336 
thiamine therapy | 120 | 336 
thiamine deficiency-associated neuropathy | 0 | 0 
GBS treatment | -720 | 120 
IVIG therapy | 0 | 120 
thiamine supplementation | 120 | 336 
neurologic symptoms | 0 | 0 
neurologic function | 192 | 336 
encephalopathy | 120 | 120 
ascending lower extremity weakness | -720 | 0 
cerebrospinal fluid (CSF) findings | 0 | 0 
intravenous immunoglobulin (IVIG) treatment | 0 | 120 
thiamine supplementation | 120 | 336 
central neurologic function | 192 | 336 
peripheral neurologic function | 192 | 336 
recovery | 192 | 336 
thiamine deficiency | -720 | 336 
beriberi | -720 | 336 
Guillain-Barré syndrome (GBS) | -720 | 120 
mimic | 0 | 0 
case reports | 0 | 0 
thiamine levels | 168 | 168 
thiamine repletion | 120 | 336 
thiamine therapy | 120 | 336 
thiamine deficiency-associated neuropathy | 0 | 0 
GBS treatment | -720 | 120 
IVIG therapy | 0 | 120 
thiamine supplementation | 120 | 336 
neurologic symptoms | 0 | 0 
neurologic function | 192 | 336 
encephalopathy | 120 | 120 
ascending lower extremity weakness | -720 | 0 
cerebrospinal fluid (CSF) findings | 0 | 0 
intravenous immunoglobulin (IVIG) treatment | 0 | 120 
thiamine supplementation | 120 | 336 
central neurologic function | 192 | 336 
peripheral neurologic function | 192 | 336 
recovery | 192 | 336 
thiamine deficiency | -720 | 336 
beriberi | -720 | 336 
Guillain-Barré syndrome (GBS) | -720 | 120 
mimic | 0 | 0 
case reports | 0 | 0 
thiamine levels | 168 | 168 
thiamine repletion | 120 | 336 
thiamine therapy | 120 | 336 
thiamine deficiency-associated neuropathy | 0 | 0 
GBS treatment | -720 | 120 
IVIG therapy | 0 | 120 
thiamine supplementation | 120 | 336 
neurologic symptoms | 0 | 0 
neurologic function | 192 | 336 
encephalopathy | 120 | 120 
ascending lower extremity weakness | -720 | 0 
cerebrospinal fluid (CSF) findings | 0 | 0 
intravenous immunoglobulin (IVIG) treatment | 0 | 120 
thiamine supplementation | 120 | 336 
central neurologic function | 192 | 336 
peripheral neurologic function | 192 | 336 
recovery | 192 | 336 
thiamine deficiency | -720 | 336 
beriberi | -720 | 336 
Guillain-Barré syndrome (GBS) | -720 | 120 
mimic | 0 | 0 
case reports | 0 | 0 
thiamine levels | 168 | 168 
thiamine repletion | 120 | 336 
thiamine therapy | 120 | 336 
thiamine deficiency-associated neuropathy | 0 | 0 
GBS treatment | -720 | 120 
IVIG therapy | 0 | 120 
thiamine supplementation | 120 | 336 
neurologic symptoms | 0 | 0 
neurologic function | 192 | 336 
encephalopathy | 120 | 120 
ascending lower extremity weakness | -720 | 0 
cerebrospinal fluid (CSF) findings | 0 | 0 
intravenous immunoglobulin (IVIG) treatment | 0 | 120 
thiamine supplementation | 120 | 336 
central neurologic function | 192 | 336 
peripheral neurologic function | 192 | 336 
recovery | 192 | 336 
thiamine deficiency | -720 | 336 
beriberi | -720 | 336 
Guillain-Barré syndrome (GBS) | -720 | 120 
mimic | 0 | 0 
case reports | 0 | 0 
thiamine levels | 168 | 168 
thiamine repletion | 120 | 336 
thiamine therapy | 120 | 336 
thiamine deficiency-associated neuropathy | 0 | 0 
GBS treatment | -720 | 120 
IVIG therapy | 0 | 120 
thiamine supplementation | 120 | 336 
neurologic symptoms | 0 | 0 
neurologic function | 192 | 336 
encephalopathy | 120 | 120 
ascending lower extremity weakness | -720 | 0 
cerebrospinal fluid (CSF) findings | 0 | 0 
intravenous immunoglobulin (IVIG) treatment | 0 | 120 
thiamine supplementation | 120 | 336 
central neurologic function | 192 | 336 
peripheral neurologic function | 192 | 336 
recovery | 192 | 336 
thiamine deficiency | -720 | 336 
beriberi | -720 | 336 
Guillain-Barré syndrome (GBS) | -720 | 120 
mimic | 0 | 0 
case reports | 0 | 0 
thiamine levels | 168 | 168 
thiamine repletion | 120 | 336 
thiamine therapy | 120 | 336 
thiamine deficiency-associated neuropathy | 0 | 0 
GBS treatment | -720 | 120 
IVIG therapy | 0 | 120 
thiamine supplementation | 120 | 336 
neurologic symptoms | 0 | 0 
neurologic function | 192 | 336 
encephalopathy | 120 | 120 
ascending lower extremity weakness