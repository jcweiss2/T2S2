73 years old | 0
male | 0
admitted to the hospital | 0
painless jaundice | -168
elevated liver functions test | -168
obstructive cholestatic pattern | -168
intrahepatic duct dilatation | 0
hypodense metastatic lesions | 0
mass effect on the common hepatic duct | 0
presumed primary cholangiocarcinoma | 0
subjective heaviness to his eyes | 0
ERCP | 24
stent insertion | 24
biliary obstruction improved | 24
cytology brushing | 24
undagnostic cytology | 24
partial ptosis of the left eyelid | 48
complete ptosis of the right eyelid | 48
binocular diplopia | 48
retro-orbital pain | 48
partial left CNIII palsy | 48
complete right CNIII palsy | 48
CT scan | 48
no intracranial lesions | 48
MRI of the brain and orbits | 72
subtle bilateral nodular lesions involving the CS | 72
18F-FDG PET/CT | 72
diffuse extensive nodal and extranodal disease | 72
multiple abdominal organs involvement | 72
bone involvement | 72
soft tissues involvement | 72
staging 18F-FDG PET/CT | 72
bilateral intense avidity of the CS | 72
targeted fine needle aspiration biopsies | 96
left level III cervical node biopsy | 96
hepatic lesion biopsy | 96
B cells with positive expression of CD10, CD19, CD20, and CD23 | 96
Ki67 proliferation index was 90% | 96
c-MYC gene rearrangement on FISH studies | 96
BL diagnosis | 96
CSF analysis | 96
negative for malignant cells | 96
hyper-CVAD chemotherapy | 120
neutropenic sepsis | 144
admission to intensive care unit | 144
de-escalation to mini R-CHOP | 168
R-CHOP | 192
intrathecal methotrexate | 192
restaging 18F-FDG PET/CT | 720
complete resolution of generalized BL deposits | 720
return to normal metabolic activity | 720
recovered full function of bilateral oculomotor nerves | 720
clinical remission | 720