23 years old | 0
male | 0
history of methicillin-resistant Staphylococcus aureus (MRSA) impetigo | -8760
right tibia fracture | -8760
intramedullary fixation (IMN) | -8760
interlocking screws removed | -840
skin irritation | -840
pain | -840
redness and swelling at the surgical site | -672
stitch abscess | -672
cultures from the surgical site were positive for MRSA | -672
oral antibiotic treatment | -672
fever | -504
right groin pain | -504
viral infection | -504
systemic fever | -336
myalgia | -336
difficult and painful ambulation | -336
right forearm cellulitis | -336
right sudden onset uveitis | -336
systemic rash | -336
right hip lymphadenopathy | -336
increased CRP | -336
elevated WBC count | -336
hepatic enzymes elevation | -336
lactic dehydrogenase (LDH) elevation | -336
creatine phosphokinase (CPK) elevation | -336
intravenous (IV) antibiotics | -336
deterioration of medical condition | -336
positron emission tomography-computed tomography (PET-CT) scan | -336
OIM abscess with systemic manifestations | -336
blood cultures were positive for MRSA bacteria | -336
hemodynamic deterioration | -336
fulminant MRSA sepsis | -336
admitted to the intensive care unit (ICU) | -336
ultrasound-guided drainage | -312
full-body CT scan | -288
enlargement of the abscesses diameter | -288
persistent fever | -288
elevated CRP level | -288
elevated WBC count | -288
surgical intervention | -264
combined approach of Smith-Peterson and modified Stoppa | -264
surgical planning | -264
general anaesthesia with muscle relaxant | -264
surgical technique | -264
Stoppa approach | -264
Smith-Peterson approach | -264
drainage and debridement of the OIM | -264
lavage for the pelvic brim | -264
improvement of general condition | -240
less frequent fever spikes | -240
decrease in CRP and WBC levels | -240
additional antibiotic treatment | -240
almost complete recovery | 0
ambulation without pain or functional limitations | 0
return to daily activities | 0