25 years old | 0
male | 0
history of intravenous drug abuse | -672
fevers | -72
back pain | -72
abdominal pain | -72
bilateral LE swelling | -72
sinus tachycardia | -72
ileofemoral and femoropopliteal acute-on-chronic deep vein thrombosis | -72
leukocytosis | -72
MRSA bacteremia | -72
tenderness to palpation in the epigastrium | -72
locally palpable thrill | -72
anasarca | -72
phlegmasia alba dolens of the bilateral LEs | -72
admitted to the hospital | 0
infrarenal MAAA | 0
spontaneous decompression via erosion into the IVC | 0
giant aortocaval fistula | 0
diminished distal arterial flow | 0
cavernous transformation of the ileofemoral venous network | 0
symmetrically diminished ankle-brachial indexes | 0
dampened aortoiliac pulse-volume recordings | 0
no evidence of active vegetation on echocardiography | 0
temporizing EVAR | 12
endovascular aneurysm repair | 12
deployment of a Gore C3 modular bifurcated endograft | 12
elimination of the aortocaval fistula | 12
immediate normalization of heart rate | 12
ascending ileofemoral venogram | 12
caval compression by the aneurysm sac | 12
multiple significant draining venous collaterals | 12
acute-on-chronic ileofemoral thrombosis | 12
refractory to catheter-directed mechanical thrombectomy | 12
open thrombectomy via common femoral venotomy and Esmarch compression | 12
hemodynamic stability achieved | 12
resolution of tachycardia | 12
phlegmasia improved | 72
leukocytosis resolved | 144
bilateral axillary unifemoral bypass grafts | 168
extra-anatomic bypass | 168
ligation of the aortic stump and the IVC | 168
explant of the temporizing endograft | 168
open repair of the mycotic aneurysm | 168
wide debridement of the MAAA | 168
surgical repair of the aortocaval fistula | 168
recovered in the intensive care unit | 192
discharged home | 240
follow-up at 1 month postoperatively | 720
follow-up at 3 months postoperatively | 2160
smooth recovery | 2160
no complications | 2160