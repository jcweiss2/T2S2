Here is the table of events and timestamps:

| Event | Timestamp |
| --- | --- |
| 18 years old | 0 |
| male | 0 |
| admitted to the hospital | 0 |
| abruptio placenta | -31 |
| emergency cesarean delivery | -31 |
| weighed 1090 g | -31 |
| Apgar values of 4 and 8 | -31 |
| hypothyroidism | -31 |
| gestational diabetes | -31 |
| group B streptococcal urine infection | -31 |
| antibiotics | -31 |
| mild respiratory distress | -1 |
| respiration rate of 65 breaths per min | -1 |
| chest retraction | -1 |
| CPAP machine | -1 |
| 6 positive end expiratory pressures and 30% inspired oxygen | -1 |
| sent to the Neonatal Intensive Care Unit (NICU) | -1 |
| cloudy eyes | 0 |
| ectropion | 0 |
| dry ichthyotic skin | 0 |
| typical male genitalia | 0 |
| bilaterally undescended testicles | 0 |
| height, weight, and head circumference | 0 |
| temperature 36.2°C | 0 |
| neurologically fine | 0 |
| heart rate 167 beats per min | 0 |
| pulsations well felt | 0 |
| CPAP with 30% FIO2 | 0 |
| breath sounds from both sides of the lung equal | 0 |
| no organomegaly in the abdomen | 0 |
| blood count, electrolytes, and liver function normal | 0 |
| respiratory distress syndrome | 0 |
| ground-glass opacity on the X-ray | 0 |
| minor respiratory acidosis | 0 |
| surfactant dosage | 0 |
| continued to receive CPAP assistance | 0 |
| bowel movement at 12 h old | 12 |
| trophic feeding | 12 |
| breast milk | 12 |
| weaned from 40% to 21% FIO2 | 12 |
| abdominal distension | 6 |
| tachycardia | 6 |
| tachypnea | 6 |
| thrombocytopenia | 6 |
| neutropenia | 6 |
| raised C-reactive protein level of 70 mg/L | 6 |
| meropenem and vancomycin | 6 |
| antibiotics escalated | 6 |
| stopped tropic feeding | 6 |
| restarted feeding at a rate of 30 mL/kg/day | 6 |
| weaned from CPAP | 14 |
| high-flow oxygen treatment | 14 |
| relapses of unexplained apnea | 21 |
| CPAP | 21 |
| FIO2 30% | 21 |
| septic examination negative | 21 |
| brain magnetic resonance imaging (MRI) normal | 21 |
| nasogastric tube | 21 |
| around half of his nutritional requirements | 21 |
| occasional breast milk and preterm formula | 21 |
| pale stools | 21 |
| neonatologist recommended a neonatal cholestasis workup | 21 |
| conjugated hyperbilirubinemia | 21 |
| total bilirubin 69.8 umol/L | 21 |
| negative septic workups | 21 |
| genetic studies on neonatal cholestasis | 21 |
| progressive familial intrahepatic cholestasis and ALGS | 21 |
| X-ray of the spine, echocardiogram, and eye test normal | 21 |
| skull X-ray revealed craniosynostosis | 21 |
| hepatosplenomegaly and signs of biliary atresia not seen | 21 |
| normal-appearing gallbladder | 21 |
| no signs of intrahepatic or extrahepatic biliary tree dilatation | 21 |
| albumin level began to decline | 21 |
| bilirubin, AST, and ALT levels rose | 21 |
| multiple albumin infusions necessary | 21 |
| ursodeoxycholic acid (30 mg/kg/day) | 21 |
| infectious etiology investigation conducted | 21 |
| results unremarkable | 21 |
| TSH, T3, T4, and cortisol levels normal | 21 |
| metabolic disorders evaluated and found to be negative | 21 |
| galactosemia and tyrosinemia type 1 | 21 |
| micropenis not detected | 21 |
| whole genomic sequence sent to a geneticist | 56 |
| caffeine and hemoglobin optimization | 56 |
| failed to manage recurrent apnea and bradycardia | 56 |
| phenobarbitone used as an empirical treatment | 56 |
| severe cyanosis, apnea, and bradycardia | 84 |
| 3 min of aggressive cardio-respiratory resuscitation | 84 |
| intubation and mechanical breathing | 84 |
| epinephrine provided | 84 |
| septic shock, multiorgan failure, and evidence of DIC | 84 |
| acute renal damage and capillary leak syndrome | 84 |
| high C-reactive protein level of 223.3 mg/L | 84 |
| died after 100 days in the hospital | 100 |
| unable to establish an etiology for the cholestatic liver illness | 100 |
| Enterobacter cloacae, gram-negative sepsis | 100 |
| diagnostic puzzle solved a week after his death | 107 |
| autosomal dominant ALGS2 caused by a pathogenic variant in the NOTCH2 gene | 107 |
| c.1076c>T (Ser359Phe) chr1: 120512166 | 107 |
| sampled blood with genomic DNA exons and intron borders | 107 |
| sequenced using the next-generation sequencing (NGS) illumina system | 107 |
| average of 80-fold coverage | 107 |
| most areas of interest covered by 15-fold coverage | 107 |
| nearly 96% covered by 20-fold coverage | 107 |
| NGS data used to align the HG19 genome assembly | 107 |
| in-house bioinformatics programs used to call and annotate genetic variants | 107 |
| detected minor alleles with less than 1% frequency in gnomAD | 107 |
| single nucleotide variants and indels checked against internal and external databases | 107 |
| automatic evidence category ratings used to classify variations | 107 |
| in-house quality score used to compare the wild-type sequence | 107 |
| variants that failed the quality score verified using PCR amplification and conventional Sanger sequencing | 107 |
| NOTCH2 gene heterozygous missense variant c.1076c>T p. (Ser359Phe) | 107 |
| results in an amino acid exchange | 107 |
| according to 8 of 10 bioinformatics in silico techniques, this variation is deleterious | 107 |
| NOTCH2 gene on chromosome 1p12 | 107 |
| responsible for Alagille syndrome 2 (ALGS2) | 107 |
| characterized by hepatic bile duct paucity and cholestasis | 107 |
| cardiac, skeletal, and ophthalmological abnormalities | 107 |
| caused by pathogenic mutations in the NOTCH2 gene | 107 |
| patients’ phenotypes seem to be dependent on the information supplied | 107 |
| ALGS2 diagnosis supported by the phenotype of patients | 107 |
| segregation study of the discovered variation in patients necessary | 107 |
| separate study of afflicted and unaffected family members beneficial | 107 |
| genetic counseling for the whole family crucial | 107 |
| Sorting Intolerant from Tolerant (SIFT) score of 0.032 | 107 |
| SIFT score interpreted as detrimental | 107 |
| Mutation Taster score of 1 | 107 |
| Combined Annotation Dependent Depletion tool score of 27.2 | 107 |
| Deep Artificial Neural Network score of 1 | 107 |
| Functional Analysis via Hidden Markov Models score of −2.63 | 107 |
| predicted pathogenic mutation for our case | 107 |
| TPN-associated cholestasis | 21 |
| direct serum bilirubin concentration of more than 34 mmol/L | 21 |
| independent of disease-related liver enzyme abnormalities | 21 |
| TPN duration, birth weight, antibiotic duration, | 21 |
| feeding, amino acids, and lipids identified as possible exposures | 21 |
| adjusted lipid infusion to 0.5 g/kg/day | 21 |
| increased carbohydrate intake to 15 kcal/kg/day | 21 |
| carnitine supplementation | 21 |
| ursodeoxycholic acid at 30 mg/kg/day | 21 |
| unable to alleviate the patient’s cholestasis | 21 |
| biliary atresia | 21 |
| symptoms such as conjugated hyperbilirubinemia | 21 |
| liver transaminases such as GGTP | 21 |
| pale stool | 21 |
| abdominal ultrasound repeated | 21 |
| gallbladder neither tiny nor nonexistent | 21 |
| normal-appearing gallbladder | 21 |
| lack of a triangular-cord sign | 21 |
| no evidence of intrahepatic or extrahepatic biliary tree dilatation | 21 |
| liver function steadily worsened | 21 |
| bilirubin, AST, and ALT levels rose | 21 |
| serum albumin fell | 21 |
| multiple albumin infusions necessary | 21 |
| ursodeoxycholic acid (30 mg/kg/day) | 21 |
| comprehensive examination found nothing wrong | 21 |
| all infectious etiologies, including TORCH and hepatitis A, B, and C | 21 |
| negative | 21 |
| TSH, T3, T4, and cortisol levels normal | 21 |
| pertinent metabolic illnesses evaluated and found to be negative | 21 |
| galactosemia and tyrosinemia type 1 | 21 |
| no anomalies observed in a thorough metabolic examination | 21 |
| blood amino acid levels, urine organic acid levels, and tandem mass spectrometry | 21 |
| normal | 21 |
| Fasting serum amino acid levels raised | 21 |
| several amino acids | 21 |
| anomalies thought to be caused by liver failure | 21 |
| investigation failed to confirm the diagnosis of panhypopituitarism | 21 |
| brain MRI normal | 21 |
| whole-exome sequencing | 56 |
| ALGS is a multisystem illness | 56 |
| affects 1 in every 30 000 babies | 56 |
| chronic cholestasis, caused by the absence of intrahepatic bile ducts | 56 |
| congenital heart disease of the pulmonary outflow tract and the vasculature | 56 |
| butterfly vertebrae | 56 |
| broad forehead | 56 |
| posterior embryotoxon and/or anterior segment abnormalities of the eyes | 56 |
| pigmentary retinopathy | 56 |
| anomalies of the basilar, carotid, and middle cerebral arteries | 56 |
| up to 15% of cases of minor head trauma-related intracranial bleeding | 56 |
| structural and functional renal defects | 56 |
| including cysts, ureteropelvic obstructions, and renal tubular acidosis | 56 |
| ALGS patients with NOTCH2 mutations and those with JAG1 mutations | 56 |
| diversity in the expression levels of the affected systems | 56 |
| liver malformations universal in NOTCH2 patients | 56 |
| ophthalmological defects and renal anomalies identical to that of JAG1 patients | 56 |
| NOTCH2 group had a tendency toward less cardiac involvement | 56 |
| 60.3% vs 100% in JAG1 | 56 |
| NOTCH2 probands showed a significantly lower degree of penetrance | 56 |
| vertebral anomalies (10%) and facial features (20%) | 56 |
| compared to the JAG1 group | 56 |
| NOTCH2 gene variants associated with Hajdu-Cheney syndrome | 56 |
| Serpentine fibula polycystic renal syndrome | 56 |
| several types of cancer | 56 |
| ALGS in our case recognized using the new ALGS genetic foundation’s diagnostic criteria | 56 |
| presence of a disease-causing mutation in the NOTCH2 gene | 56 |
| heterozygous variant c.1076c>T (Ser359Phe) chr1: 120512166 | 56 |
| 1 critical clinical characteristic of cholestasis | 56 |
| cholestasis occurs when conjugated bilirubin exceeds 1 mg/dL | 56 |
| total serum bilirubin less than 5 mg/dL | 56 |
| or when conjugated bilirubin exceeds 20% of total bilirubin over 5 mg/dL | 56 |
| total bilirubin was high (4.08 mg/dL, or 69.8 umol/L) | 56 |
| direct bilirubin was 1.27 mg/dL | 56 |
| increase of more than 20% since the start of the third week | 56 |
| NOTCH2 mutations can be difficult to diagnose | 56 |
| diversity of alterations, as well as the broad range of penetrance and clinical symptoms | 56 |
| NOTCH2 mutations may have a milder phenotype | 56 |
| compared to JAG1 mutations | 56 |
| NOTCH2 mutations may have a lower incidence of cardiac involvement | 56 |
| and vertebral malformations | 56 |
| NOTCH2 mutations may have a lower incidence of facial features | 56 |
| NOTCH2 mutations may be associated with other conditions | 56 |
| such as Hajdu-Cheney syndrome | 56 |
| Serpentine fibula polycystic renal syndrome | 56 |
| several types of cancer | 56 |
| NOTCH2 mutations may have a variable phenotype | 56 |
| depending on the specific mutation and the individual patient | 56 |
| NOTCH2 mutations may be associated with a range of clinical features | 56 |
| including liver disease, ophthalmological abnormalities, and renal defects | 56 |
| NOTCH2 mutations may be associated with a range of systemic features | 56 |
| including cardiac, skeletal, and ophthalmological abnormalities | 56 |
| NOTCH2 mutations may be associated with a range of genetic syndromes | 56 |
| including Hajdu-Cheney syndrome and Serpentine fibula polycystic renal syndrome | 56 |
| NOTCH2 mutations may be associated with an increased risk of cancer | 56 |
| NOTCH2 mutations may be associated with a range of other conditions | 56 |
| including liver disease, ophthalmological abnormalities, and renal defects | 56 |
| NOTCH2 mutations may be associated with a range of systemic features | 56 |
| including cardiac, skeletal, and ophthalmological abnormalities | 56 |
| NOTCH2 mutations may be associated with a range of genetic syndromes | 56 |
| including Hajdu-Cheney syndrome and Serpentine fibula polycystic renal syndrome | 56 |
| NOTCH2 mutations may be associated with an increased risk of cancer | 56 |
| NOTCH2 mutations may be associated with a range of other conditions | 56 |
| including liver disease, ophthalmological abnormalities, and renal defects | 56 |
| NOTCH2 mutations may be associated with a range of systemic features | 56 |
| including cardiac, skeletal, and ophthalmological abnormalities | 56 |
| NOTCH2 mutations may be associated with a range of genetic syndromes | 56 |
| including Hajdu-Cheney syndrome and Serpentine fibula polycystic renal syndrome | 56 |
| NOTCH2 mutations may be associated with an increased risk of cancer | 56 |
| NOTCH2 mutations may be associated with a range of other conditions | 56 |
| including liver disease, ophthalmological abnormalities, and renal defects | 56 |
| NOTCH2 mutations may be associated with a range of systemic features | 56 |
| including cardiac, skeletal, and ophthalmological abnormalities | 56 |
| NOTCH2 mutations may be associated with a range of genetic syndromes | 56 |
| including Hajdu-Cheney syndrome and Serpentine fibula polycystic renal syndrome | 56 |
| NOTCH2 mutations may be associated with an increased risk of cancer | 56 |
| NOTCH2 mutations may be associated with a range of other conditions | 56 |
| including liver disease, ophthalmological abnormalities, and renal defects | 56 |
| NOTCH2 mutations may be associated with a range of systemic features | 56 |
| including cardiac, skeletal, and ophthalmological abnormalities | 56 |
| NOTCH2 mutations may be associated with a range of genetic syndromes | 56 |
| including Hajdu-Cheney syndrome and Serpentine fibula polycystic renal syndrome | 56 |
| NOTCH2 mutations may be associated with an increased risk of cancer | 56 |
| NOTCH2 mutations may be associated with a range of other conditions | 56 |
| including liver disease, ophthalmological abnormalities, and renal defects | 56 |
| NOTCH2 mutations may be associated with a range of systemic features | 56 |
| including cardiac, skeletal, and ophthalmological abnormalities | 56 |
| NOTCH2 mutations may be associated with a range of genetic syndromes | 56 |
| including Hajdu-Cheney syndrome and Serpentine fibula polycystic renal syndrome | 56 |
| NOTCH2 mutations may be associated with an increased risk of cancer | 56 |
| NOTCH2 mutations may be associated with a range of other conditions | 56 |
| including liver disease, ophthalmological abnormalities, and renal defects | 56 |
| NOTCH2 mutations may be associated with a range of systemic features | 56 |
| including cardiac, skeletal, and ophthalmological abnormalities | 56 |
| NOTCH2 mutations may be associated with a range of genetic syndromes | 56 |
| including Hajdu-Cheney syndrome and Serpentine fibula polycystic renal syndrome | 56 |
| NOTCH2 mutations may be associated with an increased risk of cancer | 56 |
| NOTCH2 mutations may be associated with a range of other conditions | 56 |
| including liver disease, ophthalmological abnormalities, and renal defects | 56 |
| NOTCH2 mutations may be associated with a range of systemic features | 56 |
| including cardiac, skeletal, and ophthalmological abnormalities | 56 |
| NOTCH2 mutations may be associated with a range of genetic syndromes | 56 |
| including Hajdu-Cheney syndrome and Serpentine fibula polycystic renal syndrome | 56 |
| NOTCH2 mutations may be associated with an increased risk of cancer | 56 |
| NOTCH2 mutations may be associated with a range of other conditions | 56 |
| including liver disease, ophthalmological abnormalities, and renal defects | 56 |
| NOTCH2 mutations may be associated with a range of systemic features | 56 |
| including cardiac, skeletal, and ophthalmological abnormalities | 56 |
| NOTCH2 mutations may be associated with a range of genetic syndromes | 56 |
| including Hajdu-Cheney syndrome and Serpentine fibula polycystic renal syndrome | 56 |
| NOTCH2 mutations may be associated with an increased risk of cancer | 56 |
| NOTCH2 mutations may be associated with a range of other conditions | 56 |
| including liver disease, ophthalmological abnormalities, and renal defects | 56 |
| NOTCH2 mutations may be associated with a range of systemic features | 56 |
| including cardiac, skeletal, and ophthalmological abnormalities | 56 |
| NOTCH2 mutations may be associated with a range of genetic syndromes | 56 |
| including Hajdu-Cheney syndrome and Serpentine fibula polycystic renal syndrome | 56 |
| NOTCH2 mutations may be associated with an increased risk of cancer | 56 |
| NOTCH2 mutations may be associated with a range of other conditions | 56 |
| including liver disease, ophthalmological abnormalities, and renal defects | 56 |
| NOTCH2 mutations may be associated with a range of systemic features | 56 |
| including cardiac, skeletal, and ophthalmological abnormalities | 56 |
| NOTCH2 mutations may be associated with a range of genetic syndromes | 56 |
| including Hajdu-Cheney syndrome and Serpentine fibula polycystic renal syndrome | 56 |
| NOTCH2 mutations may be associated with an increased risk of cancer | 56 |
| NOTCH2 mutations may be associated with a range of other conditions | 56 |
| including liver disease, ophthalmological abnormalities, and renal defects | 56 |
| NOTCH2 mutations may be associated with a range of systemic features | 56 |
| including cardiac, skeletal, and ophthalmological abnormalities | 56 |
| NOTCH2 mutations may be associated with a range of genetic syndromes | 56 |
| including Hajdu-Cheney syndrome and Serpentine fibula polycystic renal syndrome | 56 |
| NOTCH2 mutations may be associated with an increased risk of cancer | 56 |
| NOTCH2 mutations may be associated with a range of other conditions | 56 |
| including liver disease, ophthalmological abnormalities, and renal defects | 56 |
| NOTCH2 mutations may be associated with a range of systemic features | 56 |
| including cardiac, skeletal, and ophthalmological abnormalities | 56 |
| NOTCH2 mutations may be associated with a range of genetic syndromes | 56 |
| including Hajdu-Cheney syndrome and Serpentine fibula polycystic renal syndrome | 56 |
| NOTCH2 mutations may be associated with an increased risk of cancer | 56 |
| NOTCH2 mutations may be associated with a range of other conditions | 56 |
| including liver disease, ophthalmological abnormalities, and renal defects | 56 |
| NOTCH2 mutations may be associated with a range of systemic features | 56 |
| including cardiac, skeletal, and ophthalmological abnormalities | 56 |
| NOTCH2 mutations may be associated with a range of genetic syndromes | 56 |
| including Hajdu-Cheney syndrome and Serpentine fibula polycystic renal syndrome | 56 |
| NOTCH2 mutations may be associated with an increased risk of cancer | 56 |
| NOTCH2 mutations may be associated with a range of other conditions | 56 |
| including liver disease, ophthalmological abnormalities, and renal defects | 56 |
| NOTCH2 mutations may be associated with a range of systemic features | 56 |
| including cardiac, skeletal, and ophthalmological abnormalities | 56 |
| NOTCH2 mutations may be associated with a range of genetic syndromes | 56 |
| including Hajdu-Cheney syndrome and Serpentine fibula polycystic renal syndrome | 56 |
| NOTCH2 mutations may be associated with an increased risk of cancer | 56 |
| NOTCH2 mutations may be associated with a range of other conditions | 56 |
| including liver disease, ophthalmological abnormalities, and renal defects | 56 |
| NOTCH2 mutations may be associated with a range of systemic features | 56 |
| including cardiac, skeletal, and ophthalmological abnormalities | 56 |
| NOTCH2 mutations may be associated with a range of genetic syndromes | 56 |
| including Hajdu-Cheney syndrome and Serpentine fibula polycystic renal syndrome | 56 |
| NOTCH2 mutations may be associated with an increased risk of cancer | 56 |
| NOTCH2 mutations may be associated with a range of other conditions | 56 |
| including liver disease, ophthalmological abnormalities, and renal defects | 56 |
| NOTCH2 mutations may be associated with a range of systemic features | 56 |
| including cardiac, skeletal, and ophthalmological abnormalities | 56 |
| NOTCH2 mutations may be associated with a range of genetic syndromes | 56 |
| including Hajdu-Cheney syndrome and Serpentine fibula polycystic renal syndrome | 56 |
| NOTCH2 mutations may be associated with an increased risk of cancer | 56 |
| NOTCH2 mutations may be associated with a range of other conditions | 56 |
| including liver disease, ophthalmological abnormalities, and renal defects | 56 |
| NOTCH2 mutations may be associated with a range of systemic features | 56 |
| including cardiac, skeletal, and ophthalmological abnormalities | 56 |
| NOTCH2 mutations may be associated with a range of genetic syndromes | 56 |
| including Hajdu-Cheney syndrome and Serpentine fibula polycystic renal syndrome | 56 |
| NOTCH2 mutations may be associated with an increased risk of cancer | 56 |
| NOTCH2 mutations may be associated with a range of other conditions | 56 |
| including liver disease, ophthalmological abnormalities, and renal defects | 56 |
| NOTCH2 mutations may be associated with a range of systemic features | 56 |
| including cardiac, skeletal, and ophthalmological abnormalities | 56 |
| NOTCH2 mutations may be associated with a range of genetic syndromes | 56 |
| including Hajdu-Cheney syndrome and Serpentine fibula polycystic renal syndrome | 56 |
| NOTCH2 mutations may be associated with an increased risk of cancer | 56 |
| NOTCH2 mutations may be associated with a range of other conditions | 56 |
| including liver disease, ophthalmological abnormalities, and renal defects | 56 |
| NOTCH2 mutations may be associated with a range of systemic features | 56 |
| including cardiac, skeletal, and ophthalmological abnormalities | 56 |
| NOTCH2 mutations may be associated with a range of genetic syndromes | 56 |
| including Hajdu-Cheney syndrome and Serpentine fibula polycystic renal syndrome | 56 |
| NOTCH2 mutations may be associated with an increased risk of cancer | 56 |
| NOTCH2 mutations may be associated with a range of other conditions | 56 |
| including liver disease, ophthalmological abnormalities, and renal defects | 56 |
| NOTCH2 mutations may be associated with a range of systemic features | 56 |
| including cardiac, skeletal, and ophthalmological abnormalities | 56 |
| NOTCH2 mutations may be associated with a range of genetic syndromes | 56 |
| including Hajdu-Cheney syndrome and Serpentine fibula polycystic renal syndrome | 56 |
| NOTCH2 mutations may be associated with an increased risk of cancer | 56 |
| NOTCH2 mutations may be associated with a range of other conditions | 56 |
| including liver disease, ophthalmological abnormalities, and renal defects | 56 |
| NOTCH2 mutations may be associated with a range of systemic features | 56 |
| including cardiac, skeletal, and ophthalmological abnormalities | 56 |
| NOTCH2 mutations may be associated with a range of genetic syndromes | 56 |
| including Hajdu-Cheney syndrome and Serpentine fibula polycystic renal syndrome | 56 |
| NOTCH2 mutations may be associated with an increased risk of cancer | 56 |
| NOTCH2 mutations may be associated with a range of other conditions | 56 |
| including liver disease, ophthalmological abnormalities, and renal defects | 56 |
| NOTCH2 mutations may be associated with a range of systemic features | 56 |
| including cardiac, skeletal, and ophthalmological abnormalities | 56 |
| NOTCH2 mutations may be associated with a range of genetic syndromes | 56 |
| including Hajdu-Cheney syndrome and Serpentine fibula polycystic renal syndrome | 56 |
| NOTCH2 mutations may be associated with an increased risk of cancer | 56 |
| NOTCH2 mutations may be associated with a range of other conditions | 56 |
| including liver disease, ophthalmological abnormalities, and renal defects | 56 |
| NOTCH2 mutations may be associated with a range of systemic features | 56 |
| including cardiac, skeletal, and ophthalmological abnormalities | 56 |
| NOTCH2 mutations may be associated with a range of genetic syndromes | 56 |
| including Hajdu-Cheney syndrome and Serpentine fibula polycystic renal syndrome | 56 |
| NOTCH2 mutations may be associated with an increased risk of cancer | 56 |
| NOTCH2 mutations may be associated with a range of other conditions | 56 |
| including liver disease, ophthalmological abnormalities, and renal defects | 56 |
| NOTCH2 mutations may be associated with a range of systemic features | 56 |
| including cardiac, skeletal, and ophthalmological abnormalities | 56 |
| NOTCH2 mutations may be associated with a range of genetic syndromes | 56 |
| including Hajdu-Cheney syndrome and Serpentine fibula polycystic renal syndrome | 56 |
| NOTCH2 mutations may be associated with an increased risk of cancer | 56 |
| NOTCH2 mutations may be associated with a range of other conditions | 56 |
| including liver disease, ophthalmological abnormalities, and renal defects | 56 |
| NOTCH2 mutations may be associated with a range of systemic features | 56 |
| including cardiac, skeletal, and ophthalmological abnormalities | 56 |
| NOTCH2 mutations may be associated with a range of genetic syndromes | 56 |
| including Hajdu-Cheney syndrome and Serpentine fibula polycystic renal syndrome | 56 |
| NOTCH2 mutations may be associated with an increased risk of cancer | 56 |
| NOTCH2 mutations may be associated with a range of other conditions | 56 |
| including liver disease, ophthalmological abnormalities, and renal defects | 56 |
| NOTCH2 mutations may be associated with a range of systemic features | 56 |
| including cardiac, skeletal, and ophthalmological abnormalities | 56 |
| NOTCH2 mutations may be associated with a range of genetic syndromes | 56 |
| including Hajdu-Cheney syndrome and Serpentine fibula polycystic renal syndrome | 56 |
| NOTCH2 mutations may be associated with an increased risk of cancer | 56 |
| NOTCH2 mutations may be associated with a range of other conditions | 56 |
| including liver disease, ophthalmological abnormalities, and renal defects | 56 |
| NOTCH2 mutations may be associated with a range of systemic features | 56 |
| including cardiac, skeletal, and ophthalmological abnormalities | 56 |
| NOTCH2 mutations may be associated with a range of genetic syndromes | 56 |
| including Hajdu-Cheney syndrome and Serpentine fibula polycystic renal syndrome | 56 |
| NOTCH2 mutations may be associated with an increased risk of cancer | 56 |
| NOTCH2 mutations may be associated with a range of other conditions | 56 |
| including liver disease, ophthalmological abnormalities, and renal defects | 56 |
| NOTCH2 mutations may be associated with a range of systemic features | 56 |
| including cardiac, skeletal, and ophthalmological abnormalities | 56 |
| NOTCH2 mutations may be associated with a range of genetic syndromes | 56 |
| including Hajdu-Cheney syndrome and Serpentine fibula polycystic renal syndrome | 56 |
| NOTCH2 mutations may be associated with an increased risk of cancer | 56 |
| NOTCH2 mutations may be associated with a range of other conditions | 56 |
| including liver disease, ophthalmological abnormalities, and renal defects | 56 |
| NOTCH2 mutations may be associated with a range of systemic features | 56 |
| including cardiac, skeletal, and ophthalmological abnormalities | 56 |
| NOTCH2 mutations may be associated with a range of genetic syndromes | 56 |
| including Hajdu-Cheney syndrome and Serpentine fibula polycystic renal syndrome | 56 |
| NOTCH2 mutations may be associated with an increased risk of cancer | 56 |
| NOTCH2 mutations may be associated with a range of other conditions | 56 |
| including liver disease, ophthalmological abnormalities, and renal defects | 56 |
| NOTCH2 mutations may be associated with a range of systemic features | 56 |
| including cardiac, skeletal, and ophthalmological abnormalities | 56 |
| NOTCH2 mutations may be associated with a range of genetic syndromes | 56 |
| including Hajdu-Cheney syndrome and Serpentine fibula polycystic renal syndrome | 56 |
| NOTCH2 mutations may be associated with an increased risk of cancer | 56 |
| NOTCH2 mutations may be associated with a range of other conditions | 56 |
| including liver disease, ophthalmological abnormalities, and renal defects | 56 |
| NOTCH2 mutations may be associated with a range of systemic features | 56 |
| including cardiac, skeletal, and ophthalmological abnormalities | 56 |
| NOTCH2 mutations may be associated with a range of genetic syndromes | 56 |
| including Hajdu-Cheney syndrome and Serpentine fibula polycystic renal syndrome | 56 |
| NOTCH2 mutations may be associated with an increased risk of cancer | 56 |
| NOTCH2 mutations may be associated with a range of other conditions | 56 |
| including liver disease, ophthalmological abnormalities, and renal defects | 56 |
| NOTCH2 mutations may be associated with a range of systemic features | 56 |
| including cardiac, skeletal, and ophthalmological abnormalities | 56 |
| NOTCH2 mutations may be associated with a range of genetic syndromes | 56 |
| including Hajdu-Cheney syndrome and Serpentine fibula polycystic renal syndrome | 56 |
| NOTCH2 mutations may be associated with an increased risk of cancer | 56 |
| NOTCH2 mutations may be associated with a range of other conditions | 56 |
| including liver disease, ophthalmological abnormalities, and renal defects | 56 |
| NOTCH2 mutations may be associated with a range of systemic features | 56 |
| including cardiac, skeletal, and ophthalmological abnormalities | 56 |
| NOTCH2 mutations may be associated with a range of genetic syndromes | 56 |
| including Hajdu-Cheney syndrome and Serpentine fibula polycystic renal syndrome | 56 |
| NOTCH2 mutations may be associated with an increased risk of cancer | 56 |
| NOTCH2 mutations may be associated with a range of other conditions | 56 |
| including liver disease, ophthalmological abnormalities, and renal defects | 56 |
| NOTCH2 mutations may be associated with a range of systemic features | 56 |
| including cardiac, skeletal, and ophthalmological abnormalities | 56 |
| NOTCH2 mutations may be associated with a range of genetic syndromes | 56 |
| including Hajdu-Cheney syndrome and Serpentine fibula polycystic renal syndrome | 56 |
| NOTCH2 mutations may be associated with an increased risk of cancer | 56 |
| NOTCH2 mutations may be associated with a range of other conditions | 56 |
| including liver disease, ophthalmological abnormalities, and renal defects | 56 |
| NOTCH2 mutations may be associated with a range of systemic features | 56 |
| including cardiac, skeletal, and ophthalmological abnormalities | 56 |
| NOTCH2 mutations may be associated with a range of genetic syndromes | 56 |
| including Hajdu-Cheney syndrome and Serpentine fibula polycystic renal syndrome | 56 |
| NOTCH2 mutations may be associated with an increased risk of cancer | 56 |
| NOTCH2 mutations may be associated with a range of other conditions | 56 |
| including liver disease, ophthalmological abnormalities, and renal defects | 56 |
| NOTCH2 mutations may be associated with a range of systemic features | 56 |
| including cardiac, skeletal, and ophthalmological abnormalities | 56 |
| NOTCH2 mutations may be associated with a range of genetic syndromes | 56 |
| including Hajdu-Cheney syndrome and Serpentine fibula polycystic renal syndrome | 56 |
| NOTCH2 mutations may be associated with an increased risk of cancer | 56 |
| NOTCH2 mutations may be associated with a range of other conditions | 56 |
| including liver disease, ophthalmological abnormalities, and renal defects | 56 |
| NOTCH2 mutations may be associated with a range of systemic features | 56 |
| including cardiac, skeletal, and ophthalmological abnormalities | 56 |
| NOTCH2 mutations may be associated with a range of genetic syndromes | 56 |
| including Hajdu-Cheney syndrome and Serpentine fibula polycystic renal syndrome | 56 |
| NOTCH2 mutations may be associated with an increased risk of cancer | 56 |
| NOTCH2 mutations may be associated with a range of other conditions | 56 |
| including liver disease, ophthalmological abnormalities, and renal defects | 56 |
| NOTCH2 mutations may be associated with a range of systemic features | 56 |
| including cardiac, skeletal, and ophthalmological abnormalities | 56 |
| NOTCH2 mutations may be associated with a range of genetic syndromes | 56 |
| including Hajdu-Cheney syndrome