64 years old | 0
female | 0
admitted to the hospital | 0
hypertension | -672
hypothyroidism | -672
tobacco use disorder | -672
takotsubo cardiomyopathy | -672
stroke | -672
acute abdominal pain | 0
nausea | -48
vomiting | -48
dry mucous membranes | 0
periumbilical abdominal tenderness | 0
temperature 36.4 °C | 0
blood pressure 65/34 mmHg | 0
heart rate 78 bpm | 0
oxygen saturation 96% | 0
hemoglobin 12.0 g/dL | 0
white blood cell count 19,890 μL | 0
lactic acid level 3.4 mmol/L | 0
creatinine level 2.65 mg/dL | 0
BUN 36 mg/dL | 0
CO2 22mEq/L | 0
voluminous non-bloody diarrhea | 2
CT of the abdomen and pelvis without contrast | 2
generalized colonic thickening | 2
moderate fluid distension of multiple loops of small bowel | 2
ascending colon | 2
transverse colon | 2
splenic flexure | 2
concern for stricture in the region of the proximal descending colon | 2
stool tests returned negative for Clostridium Difficile toxin | 2
fecal occult blood test was positive | 2
presumptive diagnosis of septic shock | 2
blood cultures were pending | 2
aggressive fluid resuscitation | 2
broad spectrum intravenous antibiotic coverage with piperacillin-tazobactam | 2
admission to the Intensive Care Unit for vasopressor support | 2
renal function improved | 48
repeat CT abdomen and pelvis was performed with IV contrast | 48
pancolonic thickening | 48
more marked involvement of the left side | 48
fecal calprotectin level of 1190 μg/mg | 48
positive fecal lactoferrin | 48
normal stool culture | 48
blood cultures growing gram variable rods | 48
inflammatory markers were markedly elevated | 48
erythrocyte sediment rate of 105 mm/h | 48
C-reactive protein level of 24 mg/dL | 48
D-dimer >20 μg/mlFEU | 48
downgraded to the general medical floor | 72
colonoscopy was performed | 72
scattered severe mucosal changes | 72
altered vascularity | 72
congestion | 72
friability | 72
granularity | 72
mucus | 72
deep ulcerations throughout the ascending, transverse, descending and sigmoid colon | 72
endoscopic biopsies confirmed pancolonic mucosal ulcerations | 72
most severe in the transverse and descending colon | 72
rectal sparing | 72
cytomegalovirus immunostaining was negative | 72
MRI angiography was negative for high grade stenosis | 72
diarrhea resolved | 72
abdominal pain, nausea and vomiting continued | 72
blood cultures returned positive for Fusobacterium Necrophorum | 168
remained on piperacillin-tazobactam | 168
consultation with colorectal surgery recommended against surgery | 168
discharged | 504
readmitted to a different hospital | 576
recurrent bloody diarrhea | 576
complicated by vancomycin-resistant Enterococcus bacteremia | 576
stabilized and discharged | 576
plan for follow up with the Gastroenterology team | 576
returned to our hospital with abdominal pain, voluminous diarrhea, and severe anemia | 672
repeat CT angiogram of the abdomen and pelvis revealed persistent diffuse colonic thickening | 672
antineutrophil cytoplasmic antibodies testing was negative | 672
persistent ischemic bowel disease | 672
surgical consultation again recommended deferring surgery | 672
monitoring for symptom improvement | 672
plan to repeat a colonoscopy shortly after discharge | 672
sought a second opinion closer to her home | 840
repeat colonoscopy performed four months after her initial presentation | 840
deep and serpentine ulcerations in a continuous and circumferential pattern | 840
involving the transverse and sigmoid colon | 840
sparing the rectum | 840
diagnosed with IBD | 840
prescribed steroids | 840
plans to transition to biologic therapy | 840
died a few months later at home | 1008