92 years old | 0
male | 0
admitted to the hospital | 0
diabetes mellitus | -672
systemic hypertension | -672
stroke | -672
general deterioration | 0
temperature of 34°C | 0
blood pressure of 70/30 mmHg | 0
pulse rate of 115 per minute | 0
respiratory rate of 22 per minute | 0
Glasgow Coma Scale of 8 out of 15 | 0
urinary tract infection | 0
septic shock | 0
intravenous fluids | 0
vasopressors | 0
mechanical ventilation | 0
imipenem-cilastatin | 0
ciprofloxacin | 0
ESBL-producing Escherichia coli | 0
ciprofloxacin replaced with gentamicin | 24
gentamicin | 24
fever up to 38.6°C | 240
hypotension | 240
peripheral blood leukocytosis | 240
dull percussion sound | 240
reduced breath sounds in the left lung | 240
left lung consolidation with a large pleural effusion | 240
pigtail catheter inserted | 240
pleural effusion drained | 240
protein at 52.0 g/L | 240
lactate dehydrogenase at 1477 IU/L | 240
pH at 7.0 | 240
white blood cells at 8450 | 240
96% neutrophils | 240
ventilator-associated pneumonia | 240
pleurisy | 240
colistin methanesulfonate | 240
imipenem-cilastatin | 240
pneumothorax | 264
pigtail catheter replaced with intercostal chest drain | 264
ESBL-producing E. coli | 264
carbapenem-resistant Acinetobacter baumannii | 264
intra-pleural colistin methanesulfonate | 336
febrile | 336
high dose vasopressor infusions | 336
lack of clinical improvement | 336
intra-pleural colistin methanesulfonate | 336
improvement in the patient’s condition | 408
peripheral white blood cell count to 8.8×10^9/L | 408
reduced need for ventilation | 408
successful discontinuation of the vasopressor support | 408
Proteus mirabilis | 408
minimum inhibitory concentrations of imipenem and meropenem | 408
switch from imipenem-cilastatin to meropenem | 408
intra-pleural and intravenous colistin methanesulfonate therapies discontinued | 448
meropenem continued | 448
culture of pleural fluid obtained on day 37 | 456
intercostal drain removed | 504
follow-up chest x-ray showed the resolution of the previously identified signs of infection and effusion | 504
acute myocardial ischemia | 1008
passed away | 1008