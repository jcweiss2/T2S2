35 years old|0
male|0
admitted to the emergency department|0
right-sided upper back pain|0
flank pain|0
cupping procedure|-24
intermittent fevers|-1008
cough|-1008
anorexia|-1008
general malaise|-1008
seen multiple naturopathic physicians|-1008
urgent care visit|-168
started on azithromycin|-168
started on doxycycline|-168
presumptive diagnosis of pneumonia|-168
improvement in febrile symptoms|-168
improvement in overall well-being|-168
blood pressure 116/75 mmHg|0
heart rate 119 beats per minute|0
respiratory rate 20 breaths per minute|0
temperature 36.2°C|0
oxygen saturation 97% on room air|0
alert|0
appropriate|0
no signs of respiratory distress|0
non-tender cupping marks on back|0
absence of breath sounds on right chest|0
soft abdomen|0
non-tender abdomen|0
chest radiograph showing 80% opacification right hemithorax|0
consistent with pneumonia|0
parapneumonic effusion|0
bedside ultrasound|0
computed tomography of chest, abdomen, pelvis|0
consultative ultrasound confirms 10.2 × 8.9 × 12.6 cm abscess in right lobe of liver|0
white blood cell count 25×109/L|0
creatinine 92 mmol/L|0
lactate 3.5 mmol/L|0
liver transaminases within normal limits|0
international normalized ratio within normal limits|0
oxygen requirements increased to 4L|0
blood pressure dropped to 90/60|0
heart rate 108|0
treated with 2 liters normal saline|0
started on levofloxacin|0
started on vancomycin|0
started on piperacillin/tazobactam|0
thoracocentesis performed|0
white blood cells 33,688 u/L with 93% neutrophils|0
initial gram stain negative|0
antibiotics switched to ceftriaxone|0
antibiotics switched to metronidazole|0
admitted to surgical intensive care unit|0
central line placement|0
interventional radiology guided liver abscess drainage|0
percutaneous drain placement|0
tube thoracostomy|0
video assisted thorascopic surgery decortication procedure|0
diaphragmatic defect found|0
continuous with hepatic abscess cavity|0
no microorganisms found on gram stain|0
no microorganisms found on subsequent cultures|0
discharged from hospital|168
intravenous ceftriaxone|168
intravenous metronidazole|168
antibiotics discontinued|672
