47 years old | 0
    woman | 0
    cirrhosis due to intestinal failure associated liver disease | 0
    referred for multivisceral transplantation | 0
    multiple small bowel resections | -1920
    visceral myopathy | -1920
    short bowel syndrome | -1920
    small intestinal bacterial overgrowth | -1920
    gastrointestinal dysmotility | -1920
    liver biopsy | -960
    advanced cirrhosis | -960
    multivisceral transplantation indicated | -960
    donor cytomegalovirus IgG negative | 0
    recipient cytomegalovirus IgG negative | 0
    methylprednisolone induction immunosuppression | 0
    alemtuzumab induction immunosuppression | 0
    prednisolone maintenance immunosuppression | 0
    tacrolimus maintenance immunosuppression | 0
    cyclosporine replacement due to posterior reversible encephalopathy syndrome | 960
    meropenem prophylaxis | 0
    vancomycin prophylaxis | 0
    liposomal amphotericin B prophylaxis | 0
    co-trimoxazole prophylaxis | 0
    acyclovir prophylaxis | 0
    Candida glabrata isolated from blood cultures | 72
    Candida glabrata isolated from drain fluid | 72
    increased liposomal amphotericin B dose | 72
    voriconazole started due to cutaneous drug reaction | 72
    prolonged period of pyrexia | 72
    intermittent bacteremia | 72
    enterococci bacteremia | 72
    Elizabethkingia meningoseptica bacteremia | 72
    Staphylococcus haemolyticus bacteremia | 72
    Escherichia coli bacteremia | 72
    voriconazole switched to micafungin | 2304
    low serum voriconazole levels | 2304
    micafungin dose increased | 2304
    diffuse maculopapular rash | 1896
    skin biopsy demonstrated graft-versus-host disease | 1896
    donor-positive lymphocytes | 1896
    rapid bone marrow failure | 2160
    frequent transfusions | 2160
    acellular bone marrow | 2160
    increased immunosuppression | 2160
    basiliximab added | 2160
    alemtuzumab added | 2160
    immunosuppression withdrawn | 2880
    haplo-identical bone marrow transplant planned | 4032
    granulocyte infusion given | 3936
    platelet increment | 3936
    dysarthria | 3936
    unilateral upper motor neurone facial nerve palsy | 3936
    cranial CT scan | 3936
    acute frontal infarct | 3936
    deterioration | 3936
    transfer to ICU | 3936
    repeat CT showing extensive infarcts | 3936
    cerebral infarct extension | 3936
    hemorrhagic transformation | 3936
    edema | 3936
    midline shift | 3936
    treatment withdrawal | 3936
    death | 3936
    invasive mucormycosis | 3936
    vasculature involvement | 3936
    parenchyma involvement | 3936
    left ventricular fungal thrombus | 3936
    micafungin received for 69 days | 0
    no time without antifungal coverage | 0
    early Candida isolates | 72
    negative fungal cultures | 0
    negative serum galactomannan levels | 0
    <|eot_id|>
    47 years old | 0
    woman | 0
    cirrhosis due to intestinal failure associated liver disease | 0
    referred for multivisceral transplantation | 0
    multiple small bowel resections | -1920
    visceral myopathy | -1920
    short bowel syndrome | -1920
    small intestinal bacterial overgrowth | -1920
    gastrointestinal dysmotility | -1920
    liver biopsy | -960
    advanced cirrhosis | -960
    multivisceral transplantation indicated | -960
    donor cytomegalovirus IgG negative | 0
    recipient cytomegalovirus IgG negative | 0
    methylprednisolone induction immunosuppression | 0
    alemtuzumab induction immunosuppression |# hello-world
Testing
Hi, I am a new to coding but i love learning new things. 
