60 years old | 0
male | 0
diabetes mellitus | 0
hypertension | 0
admitted to the hospital | 0
transurethral re-section of the prostate | 0
refractory urine retention | 0
no loin pain | 0
no fever | 0
no rigors | 0
no previous surgery | 0
no renal angle tenderness | 0
benign digital rectal examination | 0
persistent pus cells | -24
positive pansensitive Escherichia coli | -24
urethral catheter exchange | -24
levofloxacin | -24
enlarged prostate | -24
46 gm prostate | -24
transurethral resection of the prostate | 0
piperacillin/tazobactam | 0
antibiotic coverage | 0
recurrent high-grade fever | 24
left loin pain | 24
elevated septic parameters | 24
urine culture positive for Candida albicans | 24
blood culture positive for Candida albicans | 24
intravenous fluconazole | 24
no response to fluconazole | 48
CT urography | 48
left hydronephrosis | 48
filling defect in the left renal pelvis | 48
no enhancement | 48
contrast outlining the lesion | 48
suspected renal fungal ball | 48
left percutaneous nephrostomy | 72
nephrostogram | 72
filling defects in the renal pelvis | 72
whitish debris | 72
cultures from nephrostomy positive for Candida albicans | 72
cultures from urethral catheter positive for Candida albicans | 72
cultures from blood positive for Candida albicans | 72
anidulafungin | 96
100 mg anidulafungin | 96
once daily anidulafungin | 96
improved patient condition | 120
repeated blood culture negative | 120
urine from bladder positive for candida | 120
urine from nephrostomy positive for candida | 120
instillation of fluconazole | 120
300 mg fluconazole | 120
500 mL normal saline | 120
12 hours | 120
40 mL/hour | 120
7 days | 168
urine culture from nephrostomy tube no growth | 168
midstream urine mixed growth with some candida | 168
follow-up renal ultrasound | 168
normal left kidney | 168
no lesion in the pelvicalyceal system | 168
nephrostomy tube in place | 168
nephrostomy tube removed | 216
urine culture no candida growth | 216