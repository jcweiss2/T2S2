39 years old | 0
female | 0
SLE | -8760
anti-nuclear antibody | -8760
anti-Smith positive | -8760
dsDNA+ | -8760
hypocomplementemia | -8760
history of proteinuria | -8760
immune thrombocytopenic purpura | -8760
fatigue | -36
abdominal pain | -36
severely thrombocytopenic | -36
platelets 5 × 10^9/L | -36
multiple platelet transfusions | -36
IV methylprednisolone | -36
IV immunoglobulin | -36
splenectomy | -36
intra-abdominal hematoma | -36
ischemic left foot | -36
below-the-knee amputation | -36
SLE exacerbation | -36
enterocolitis | -36
sepsis | -36
transferred to intensive care unit | -36
sloughing | -24
profound hypotension | -24
transferred to hospital | 0
temperature 31.5°C | 0
heart rate 87 | 0
blood pressure 90 to 100/40 to 50 mm Hg | 0
blood oxygen saturation 99% | 0
confluent dusky Nikolsky-positive plaques | 0
denudation | 0
crusted erosions on lips | 0
crust on conjunctiva | 0
greater than 90% total body surface area denuded or Nikolsky positive | 0
severe lactic acidosis | 0
anemia | 0
hemoglobin 5.3 g/dL | 0
thrombocytopenia | 0
platelets 42 × 10^9/L | 0
coagulopathic | 0
international normalized ratio 1.3 | 0
prothrombin time 15.1 | 0
partial thromboplastin time 60.5 | 0
protein S level decreased | 0
right femoral vein deep venous thrombosis | 0
multifocal renal cortical infarctions | 0
IV methylprednisolone | 0
continuous renal replacement therapy | 0
mitral valve thickening | 0
ciprofloxacin | 0
gentamycin | 0
vancomycin | 0
prophylactic heparin | 0
biopsy of right shin | 12
full-thickness epidermal necrosis | 12
microvascular thrombi | 12
resolving interface dermatitis | 12
plasma exchange | 24
IVIg | 24
mycophenolate mofetil | 24
anticardiolipin negative | 24
anti-β2 glycoprotein I negative | 24
antiphosphatidylserine negative | 24
fever | 48
ventilator-associated pneumonia | 48
vancomycin-resistant Enterococcus bacteremia | 72
withdraw life-sustaining therapies | 96
refractory hypotension | 120
toxic epidermal necrolysis | 120
acute hemorrhagic pancreatitis | 120
extensive necrosis | 120
fat necrosis | 120