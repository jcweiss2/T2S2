52 years old | 0 | 0 
female | 0 | 0 
admitted to the hospital | 0 | 0 
abdominal pain | -48 | 0 
nausea | -48 | 0 
vomiting | -48 | 0 
increased level of liver enzyme alanine aminotransferase | -840 | -840 
positive autoimmune antibody | -840 | -840 
elevated immunoglobulin G | -840 | -840 
coarse liver surface | -840 | -840 
liver biopsy | -840 | -840 
diagnosed with overlap syndrome | -840 | -840 
started to take ursodeoxycholic acid | -840 | -728 
started to take prednisolone | -840 | -728 
reduced prednisolone | -728 | -728 
maintained ursodeoxycholic acid | -728 | 0 
maintained azathioprine | -600 | 0 
mild heartburn | -48 | -48 
abdominal pain worsened | -24 | -24 
nausea worsened | -24 | -24 
vomiting worsened | -24 | -24 
diarrhea | -24 | -24 
visited emergency room | 0 | 0 
blood pressure normal | 0 | 0 
mild fever | 0 | 0 
tachycardia | 0 | 0 
tachypnea | 0 | 0 
abdominal tenderness | 0 | 0 
reduced white blood cells | 0 | 0 
reduced platelets | 0 | 0 
decreased neutrophil level | 0 | 0 
elevated C-reactive protein level | 0 | 0 
elevated aspartate aminotransferase | 0 | 0 
elevated ALT | 0 | 0 
elevated gamma glutamyl transferase | 0 | 0 
prothrombin time international normalized ratio | 0 | 0 
contrast-enhanced abdominal CT | 0 | 0 
huge stomach with layered wall thickening | 0 | 0 
air in the stomach wall | 0 | 0 
decrease of mucosal enhancement | 0 | 0 
diagnosed with necrotizing gastritis | 0 | 0 
diagnosed with septic shock | 0 | 0 
intravenous hydration | 0.5 | 2 
antibiotic treatment | 0.5 | 2 
transferred to intensive care unit | 0.5 | 2 
inotropics | 2 | 2 
fluid treatment | 2 | 2 
heart rate slowed | 3 | 3 
bedside echocardiography | 3 | 3 
severe stress-induced cardiomyopathy | 3 | 3 
extracorporeal membrane oxygenation | 3 | 3 
cardiac arrest | 3 | 3 
cardiopulmonary resuscitation | 3 | 3 
died | 3 | 3 
necrotizing gastritis | 0 | 3 
septic shock | 0 | 3 
azathioprine side effects | -600 | 0 
steroid side effects | -840 | 0 
leukopenia | 0 | 0 
infection | 0 | 0 
abdominal pain | -48 | 0 
nausea | -48 | 0 
vomiting | -48 | 0 
diarrhea | -24 | -24 
gastrointestinal symptoms | -48 | 0 
immunosuppressant treatment | -840 | 0 
liver function tests | -840 | 0 
blood sugar | -840 | 0 
complete blood count test | -840 | 0 
liver biopsy results | -840 | -840 
overlap syndrome diagnosis | -840 | -840 
ursodeoxycholic acid treatment | -840 | -728 
prednisolone treatment | -840 | -728 
azathioprine treatment | -600 | 0 
abdominal CT results | 0 | 0 
necrotizing gastritis diagnosis | 0 | 0 
septic shock diagnosis | 0 | 0 
intravenous antibiotics | 0.5 | 2 
fluid treatment | 0.5 | 2 
inotropics treatment | 2 | 2 
extracorporeal membrane oxygenation treatment | 3 | 3 
cardiopulmonary resuscitation | 3 | 3 
death | 3 | 3