18 years old | 0
male | 0
history of mucosal resection for early gastric cancer | -672
history of partial resection for left lung cancer | -672
history of conventional drugs | -672
67 years old | 0
knee-high wild grass from a riverbed for 10 days | -720
systemic pain and fatigue | -720
fever | -720
chills | -720
watery diarrhea | -720
loss of appetite | -720
mildly disturbed consciousness | -720
decreased white blood cells (WBC) | -720
platelet counts | -720
elevated hepatic enzyme levels | -720
hemophagocytosis | -720
suspected sepsis and febrile neutropenia (FN) | -720
administered antibiotics | -720
elevated ferritin levels | -144
screened for cytomegalovirus and Epstein-Barr virus (EBV) | -144
negative blood culture | -144
bone marrow biopsy | -144
hemophagocytosis with fewer mature myeloid series cells | -144
CD3- and CD4-positive T cells | -144
MUM-1-positive lymphoid cells | -144
CD68, CD163-positive histiomonocytes | -144
diagnosed with HLH | -144
administered prednisolone (PSL) | -144
chest pain | -144
shivering | -144
fever of 39.2°C | -144
blood pressure at 88/52 mmHg | -144
HR at 89/min | -144
RR at 24/min | -144
SPO2 at 94% | -144
elevated CK levels | -144
LDH at 1,405 U/L | -144
high-sensitivity troponin I (TnI) at 271 pg/mL | -144
severe left ventricular dysfunction | -144
ST elevation in the V1-2 leads | -144
suspected SFTS | -144
RT-PCR analysis of the submitted serum detected 1.77×106 SFTSV RNA copies/mL | -144
negative-pressure room | -144
steroid pulse therapy for HLH with SFTS | -144
withdrawn from circulatory agonist and ventilator management | -168
ECG showed improvement of ST elevation in the V1-2 leads | -168
re-submitted his serum and confirmed negativity for viremia | -168
released from quarantine | -168
CAG and EMB | -168
no coronary artery stenosis was observed on CAG | -168
pathological evaluation of the EMB specimen revealed that the myocardium was mildly hypertrophic | -168
mild myofibrillar loss and disarrangement | -168
active mononuclear cell infiltration adjacent to the damaged myocardium was not observed | -168
CD3-positive T cells | -168
CD68-positive macrophages | -168
tenascin-C expression in the stroma | -168
discharged | -168
follow-up visit 1 month after discharge | -168
transthoracic echocardiography showed a slight improvement with an EF of 52.5% | -168
no heart failure | -168
admitted to the hospital | 0
admitted to the ICU | 0
administered inotropic agents and water balance management | 0
suspected sepsis and febrile neutropenia (FN) | 0
administered antibiotics | 0
suspected SFTS | 0
RT-PCR analysis of the submitted serum detected 1.77×106 SFTSV RNA copies/mL | 0
negative-pressure room | 0
steroid pulse therapy for HLH with SFTS | 0
withdrawn from circulatory agonist and ventilator management | 0
ECG showed improvement of ST elevation in the V1-2 leads | 0
re-submitted his serum and confirmed negativity for viremia | 0
released from quarantine | 0
CAG and EMB | 24
no coronary artery stenosis was observed on CAG | 24
pathological evaluation of the EMB specimen revealed that the myocardium was mildly hypertrophic | 24
mild myofibrillar loss and disarrangement | 24
active mononuclear cell infiltration adjacent to the damaged myocardium was not observed | 24
CD3-positive T cells | 24
CD68-positive macrophages | 24
tenascin-C expression in the stroma | 24
discharged | 24
follow-up visit 1 month after discharge | 24
transthoracic echocardiography showed a slight improvement with an EF of 52.5% | 24
no heart failure | 24
SFTS | -720
HLH | -720
myocarditis | -144
febrile neutropenia (FN) | -720
hemophagocytosis | -720
sepsis | -720
disseminated intravascular coagulation | -144
acute myocarditis | -144
cardiogenic shock | -144
myocardial inflammation | 24
myocardial hypertrophy | 24
myofibrillar loss and disarrangement | 24
CD3-positive T cells | 24
CD68-positive macrophages | 24
tenascin-C expression in the stroma | 24