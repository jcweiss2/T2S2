70 years old | 0
    woman | 0
    admitted to Plastic Surgery department | -24
    fever | -24
    dizziness | -24
    unstable angina | -10800
    diabetes mellitus | -10800
    third-degree burn to the sacral area | -2520
    skin flap operation | -2520
    sore at sacral area | -1440
    osteomyelitis | -1440
    pale | 0
    febrile | 0
    temperature of 38.2℃ | 0
    intermittent fever of 37.3-38.1℃ | 0
    blood pressure 110/80 mmHg | 0
    pulse 78/min | 0
    respiratory rate 20/min | 0
    peripheral WBC count 8,730/µL | 0
    hemoglobin level 8.6 g/dL | 0
    platelet count 261,000/µL | 0
    AST 7 U/L | 0
    ALT 11 U/L | 0
    alkaline phosphatase 77 U/L | 0
    blood urea nitrogen 23.4 mg/dL | 0
    creatinine 1.42 mg/dL | 0
    total protein 5.6 g/dL | 0
    albumin 2.9 g/dL | 0
    erythrocyte sedimentation rate 53 mm/hr | 0
    C-reactive protein 220.03 mg/L | 0
    urine yellow | 0
    urine turbid | 0
    positive WBC (3+) in urine | 0
    positive protein (1+) in urine | 0
    microscopic examination >60 WBCs | 0
    yeast organisms in urine | 0
    chest radiograph right pleural thickening | 0
    chest radiograph collapse of the right lower lung | 0
    abdomen and pelvic CT cystitis | 0
    abdomen and pelvic CT fluid collection | 0
    blood culture negative | 120
    urine culture Candida albicans | 0
    fever 38.1℃ on HD 32 | 768
    blood culture negative | 768
    multidrug-resistant K. pneumoniae isolated from urine | 768
    Vitek2 GN species identification | 768
    AST-N044 antimicrobial susceptibility test | 768
    resistant to most antibiotics | 768
    gentamicin susceptible | 768
    tigecycline MIC 1 µg/mL | 768
    colistin MIC 0.25 µg/mL | 768
    modified Hodge test positive | 768
    AmpC test negative | 768
    ESBL test negative | 768
    carbapenemase inhibition test APB positive | 768
    PCR blaKPC-2 gene detected | 768
    MLST ST258 | 768
    initial treatment with ertapenem | 768
    tigecycline administered | 768
    pyuria not subsided | 768
    wound not subsided | 768
    repeated isolation of MDR K. pneumoniae | 768
    treatment with colistin | 768
    clinical improvement not observed | 768
    kidney function declining | 768
    managed in ICU | 768
    expired | 2160
    septic shock | 2160
    multiorgan failure | 2160
    