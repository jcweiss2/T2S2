54 years old | 0
man | 0
chronic cough | 0
squamous cell carcinoma | 0
left lower lobe | 0
ostium secundum atrial septal defect | 0
gastroesophageal reflux disease | 0
pulmonary left lower sleeve lobectomy | 0
general anesthesia | 0
isolated lung | 0
SpO2 96%–100% | 0
monitored left radial arterial pressure | 0
monitored central venous pressure | 0
video-assisted thoracoscopy | 0
mobilized left lower lobar pulmonary artery | 0
mobilized inferior pulmonary vein division | 0
stapled left lower lobar pulmonary artery | 0
stapled inferior pulmonary vein division | 0
calcified nodules | 0
converted to open thoracotomy | 0
dissected seventh subcarinal lymph node | 0
removed entire lower left pulmonary lobe | 0
extubated | 0
spontaneous respiration | 0
arrival in PACU | 0
conscious | 0
breathing spontaneously | 0
SpO2 90% | 0
blood pressure 136/107 mmHg | 0
blood pressure dropped to 65/49 mmHg | 5
dyspneic | 5
dopamine infusion | 5
rapid fluid infusion | 5
notified thoracic surgeons | 5
blood pressure decreased to 48/37 mmHg | 10
elevated leg | 10
inferolateral ST depression | 10
jugular vein engorgement | 10
blood pressure increased to 92/71 mmHg | 30
phenylephrine injection | 30
dopamine infusion increased | 30
SpO2 decreased to 85% | 30
SpO2 increased to 93% | 30
continuous positive airway pressure | 30
blood pressure dropped to 63/51 mmHg | 105
refractory to epinephrine | 105
refractory to fluid bolus | 105
dyspnea worsening | 105
tachypnea worsening | 105
intubated | 120
chest X-ray haziness | 120
enlarged heart | 120
straightened left cardiac border | 120
jugular vein distended | 120
suspected cardiac tamponade | 120
performed TEE | 155
detected pericardial effusion | 155
attempted pericardiocentesis | 180
insufficient pericardial drainage | 180
emergency pericardial window operation | 180
suctioned pericardial fluid | 180
hemodynamics improved | 180
blood pressure 120/70 mmHg | 180
SpO2 100% | 180
no origin found | 180
recovered well | *
outpatient chest X-rays clear | *
removed entire lower left pulmonary lobe |%0
