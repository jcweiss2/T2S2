56 years old | 0
woman | 0
history of left hydronephrosis | -2928
ureteroscopy for left ureter | -2928
laparoscopy for lysis of adhesion around left ureter | -2928
abdominal discomfort | -48
abdominal distension | -48
oliguria | -48
irritable | -48
body temperature of 39.4°C | -48
pulse rate at 114 beats per minute | -48
blood pressure declined to 86/59 mm Hg | -48
respiratory rate at 28 breaths per minute | -48
oxygen saturation of 89% under oxygen inhalation | -48
no positive signs on abdominal examination | -48
white blood cell count of 15.4 × 109/L | -48
95% neutrophils | -48
5% lymphocytes | -48
platelet count of 33 × 109/L | -48
blood lactate level of 3.6 mmol/L | -48
base excess of −11.4 | -48
serum creatinine increased to 365.7 μmol/L | -48
ALT increased to 224U/L | -48
AST increased to 858U/L | -48
prothrombin time extended to 24.2 seconds | -48
C-reactive protein of 180.3 mg/L | -48
procalcitonin of 49.17 ng/mL | -48
qSOFA score of 3 points | -48
admitted to the ICU | 0
APACHE II score of 32 | 0
SOFA score of 17 | 0
diagnosis of sepsis | 0
primaxin (imipenem/cilastatin) | 0
norepinephrine | 0
hydrocortisone | 0
supplemental fluids | 0
continuous renal replacement therapy | 0
acute kidney injury (stage 3) | 0
respiratory distress | 0
oxygenation index of 184 mm Hg | 0
endotracheal intubation | 0
mechanical ventilation | 0
white blood cell count peaked at 45.3 × 109/L | 48
91.5% neutrophils | 48
1.8% lymphocytes | 48
blood culture negative | 48
urine culture negative | 48
abdominal drainage fluid culture negative | 48
vital signs improved | 48
clinical condition improved | 48
total bilirubin rose to 245.5 μmol/L | 120
direct bilirubin rose to 196.6 μmol/L | 120
liver function failure | 120
gallbladder wall edema | 120
hepatoprotective drugs | 0
supportive therapies | 0
plasma exchange | 120
plasma exchange on 4 consecutive days | 120
mechanical ventilation stopped | 216
endotracheal tube withdrawn | 216
hemodialysis treatment continued | 216
transferred back to urology department | 288
ALT of 23 U/L | 288
AST of 39 U/L | 288
TB of 99.4 μmol/L | 288
DB of 69.8 μmol/L | 288
liver function returned to normal | 360
