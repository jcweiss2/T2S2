58 years old | 0  
    male | 0  
    admitted to the hospital | 0  
    hyperpyrexia | -168  
    dyspnoea | -48  
    cough | -48  
    phlegm with blood | -48  
    hypertension | -17520  
    poultry-related exposure | -168  
    community-acquired pneumonia | -168  
    antibacterial therapy | -168  
    increased C-reactive protein | 0  
    increased procalcitonin | 0  
    leukopenia | 0  
    lymphopenia | 0  
    decreased CD3 T cells | 0  
    decreased CD4 T cells | 0  
    decreased CD8 T cells | 0  
    HIV antibody negative | 0  
    mechanical ventilation | 0  
    moxifloxacin | 0  
    cefoperazone-sulbactam | 0  
    corticosteroids | 0  
    continuous renal replacement therapy | 0  
    influenza A (H7N9) virus positive | 0  
    oseltamivir | 0  
    Staphylococcus haemolyticus bloodstream infection | 168  
    vancomycin | 168  
    imipenem/cilastatin | 168  
    caspofungin | 168  
    Pseudomonas aeruginosa | 168  
    subcutaneous emphysema | 240  
    mediastinal emphysema | 240  
    ventilator parameters decreased | 240  
    Cryptococcus neoformans positive | 384  
    cryptococcal capsular polysaccharide antigen positive | 384  
    flucytosine | 384  
    fluconazole | 384  
    voriconazole | 384  
    amphotericin B | 384  
    itraconazole | 384  
    Stenotrophomonas maltophilia positive | 936  
    septic shock | 1128  
    disseminated intravascular coagulation | 1128  
    multi-organ failure | 1128  
    death | 1128  
