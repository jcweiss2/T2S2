29 years old | 0 | 0 
male | 0 | 0 
admitted to the hospital | 0 | 0 
muscle pain | -144 | 0 
joint pain | -144 | 0 
general weakness | -144 | 0 
fever | -144 | 0 
liver dysfunction | -144 | 0 
total bilirubin 5.7 mg/dl | -144 | 0 
serum glutamic oxaloacetic transaminase 633 U/L | -144 | 0 
serum glutamic pyruvate transaminase 412 U/L | -144 | 0 
gamma-glutamyl transferase 161 U/L | -144 | 0 
lactate dehydrogenase 1668 U/L | -144 | 0 
C-reactive protein 519 mg/l | -144 | 0 
procalcitonin 1.28 ng/ml | -144 | 0 
leukocyte levels 14.8 × 10³/μl | -144 | 0 
acute respiratory failure | 0 | 0 
altered state of consciousness | 0 | 0 
continuous sedation | 0 | 336 
muscle relaxation | 0 | 336 
intubation | 0 | 336 
mechanical ventilation | 0 | 336 
FiO2 100% | 0 | 336 
SpO2 88.7% | 0 | 336 
hemodynamic instability | 0 | 168 
norepinephrine | 0 | 168 
vasopressin | 0 | 0 
broad-spectrum empirical antimicrobial therapy | 0 | 168 
meropenem | 0 | 168 
azithromycin | 0 | 168 
oseltamivir | 0 | 168 
methylprednisolone | 0 | 168 
stress ulcer prophylaxis | 0 | 168 
thromboprophylaxis | 0 | 168 
prone position | 0 | 24 
chest CT | 0 | 24 
bedside focus ultrasound | 0 | 168 
acute renal failure | 144 | 144 
CRRT | 144 | 336 
CytoSorb adsorber | 168 | 192 
septic episode | 240 | 240 
second CytoSorb therapy | 240 | 264 
norepinephrine discontinued | 192 | 192 
inflammatory marker levels decreased | 168 | 336 
CRP decreased | 168 | 336 
leukocyte levels normalized | 168 | 336 
ICU delirium | 168 | 336 
antipsychotics | 168 | 336 
percutaneous tracheostomy | 168 | 336 
ventilator weaning | 336 | 336 
discharged from MICU | 336 | 336 
transferred to general ward | 336 | 336 
transferred to rehabilitation clinic | 336 | 336 
influenza A (H1N1) | -144 | 0 
bilateral pneumonia | -144 | 0 
massive bilateral pneumonia | 0 | 0 
minimal pleural effusions | 0 | 0 
lung-protective ventilation | 0 | 336 
lung function improvement | 168 | 336 
ventilation parameters improvement | 168 | 336 
hemodynamic stabilization | 168 | 336 
inflammation control | 168 | 336 
vasopressors discontinued | 192 | 192 
inflammation markers decrease | 168 | 336 
gradual improvement | 168 | 336 
recovery | 336 | 336