90 years old | 0
male | 0
severe abdominal pain | 0
nausea | 0
vomiting | 0
inability to defecate | 0
inability to pass gas | 0
admitted to separate healthcare facilities with abdominal pain | -43200
admitted to separate healthcare facilities with constipation | -43200
no pathology found by tests and examinations | -43200
lost 5-6 kg | -8760
hypertension | 0
salt-free diet | 0
cachectic general appearance | 0
distended abdomen | 0
dry mucosae | 0
blood pressure 90/50 mmHg | 0
pulse rate 95 bpm | 0
body temperature 37.9°C | 0
marked rebound tenderness | 0
guarding in all quadrants | 0
WBC 8.890 (neutrophil: 86.1%) | 0
Hemoglobin 14 gr/dL | 0
BUN 38 mg/dL | 0
creatinine 0.8 mg/dL | 0
diffuse air-fluid levels on upright plain abdominal X-Ray | 0
physical examination findings consistent with tumoral obstruction | 0
physical examination findings consistent with viscus perforation | 0
laparotomy via midline incision | 0
abdominal exploration revealing encapsulation of all intestinal segments | 0
dense, plate-like fibrous membrane encasing whole small intestine | 0
dense adhesions between intestinal loops | 0
loop ileostomy established | 0
admitted to intensive care unit | 0
poor general status | 0
aggressive fluid replacement | 0
electrolyte replacement |8 0
administration of wide-spectrum antibiotics | 0
septic shock | 72
multiorgan failure | 72
WBC 1880/µL | 72
BUN 123 mg/dL | 72
creatinine 2.92 mg/dL | 72
albumin 2.4 gr/dL | 72
death | 72
