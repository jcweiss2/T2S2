41 years old | 0
African-American | 0
female | 0
type 2 diabetes mellitus | -672
fever | -2
nausea | -2
vomiting | -2
diarrhea | -2
mild upper-respiratory tract infection | -168
marijuana use | -168
exposed to son with flu-like symptoms | -168
no recent travel outside the United States | 0
blood pressure 115/64 mmHg | 0
heart rate 127 beats/min | 0
respiratory rate 28 breaths/min | 0
fever of 38.8°C | 0
oxygen saturation of 97% on room air | 0
weight 79 kg | 0
BMI of 32 | 0
drowsiness | 0
mild epigastric tenderness | 0
bilateral lung infiltrates | 0
sepsis | 0
disseminated intravascular coagulopathy | 0
multi-organ failure | 0
metronidazole 500 mg/IV q8h | 0
ciprofloxacin 400 mg/IV q12h | 0
progressive respiratory failure | 12
intubation | 12
acute respiratory distress syndrome | 168
anuric | 72
hemodialysis | 72
acute liver failure | 72
acute pancreatitis without necrosis | 72
multiple transfusions | 72
anemia | 72
thrombocytopenia | 72
dry-foot gangrene | 72
amputation above the toes | 72
borderline hypotension | 72
no vasopressor support | 72
pan-sensitive Streptococcus pneumoniae in blood cultures | 0
broad-spectrum antibiotics | 0
limited clinical improvement | 168
bicytopenia | 168
hypertriglyceridemia | 168
low fibrinogen | 168
hyperferritinemia | 168
intravenous immunoglobulin 100 g/IV q24h | 168
high-dose dexamethasone therapy 20 mg/IV q24h | 168
elevated sIL2 assay | 192
deferred etoposide-based regimen | 240
extubation | 240
transfer to sub-acute rehab facility | 240
critical illness-induced myopathy | 240
physical therapy | 240