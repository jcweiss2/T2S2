58 years old | 0
male | 0
admitted to the hospital | 0
high grade fever | -336
chills | -336
bilateral loin pain | -336
pain related to the left thigh | -168
diabetes mellitus | 0
history of recurrent UTI | 0
no history of stone disease | 0
creatinine 917 μmol/L | 0
hemoglobin 6.5 g/dL | 0
total leucocytic count 40.7 × 10^3 | 0
INR 1.8 | 0
creatinine kinase 447 | 0
random blood sugar 8.45 mmol/L | 0
E. coli in urine culture | 0
no growth of organisms in blood culture | 0
bilateral emphysematous pyelonephritis | 0
right kidney marked hydronephrosis | 0
multiple air locules in right kidney | 0
right ileopsoas muscle infiltration | 0
left kidney small in size | 0
multiple renal stones in left kidney | 0
multiple air locules in left kidney | 0
empirical antibiotics | 0
ICU admission | 0
broad spectrum antibiotics | 24
bilateral nephrostomy tubes fixation | 24
retroperitoneal drains | 24
clinical improvement | 48
total leucocytic count 16.6 | 48
creatinine 663 μmol/L | 48
HGB 8.2 g/dL | 48
follow up CT | 48
resolution of EP and psoas abscess | 48
general condition deteriorated | 72
retransferred to ICU | 72
profuse rectal bleeding | 72
colonoscopy | 72
patchy oozing bleeding colonic mucosa | 72
inotropes | 72
passed away | 168