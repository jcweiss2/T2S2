39 years old | 0
male | 0
admitted to hospital | 0
ingestion of drain cleaner liquid | -5
sodium hydroxide ingestion | -5
potassium hydroxide ingestion | -5
carbonyl diamide ingestion | -5
endotracheally intubated | -5
edematous oral mucosa | 0
chemical injuries to face | 0
white blood cell count of 12.9 × 10^3/μL | 0
D-dimer > 5250 ng/mL | 0
thickening and submucosal edema of esophageal and gastric wall | 0
trace para-esophageal and peri-gastric stranding and fluid | 0
no free air | 0
tracheostomy | 13
jejunostomy tube | 13
coughing during sedation-awakening trials | 13
reduction in sedatives | 13
acutely hypoxic | 18
oxygen saturation decreased to 50% | 18
pulseless electrical arrest | 18
advanced cardiopulmonary resuscitation | 18
recovery of spontaneous circulation | 18
copious amounts of frothy, yellow-tinted secretions | 18
no oral secretions | 18
nasogastric tube placement | 18
gastric cavity decompression | 18
approximately 400-500 mL of fluid suctioned | 18
esophageal stent placement | 22
acute respiratory distress syndrome | 22
recurrent septic shock | 22
aspiration pneumonia | 22
liberated from mechanical ventilation | 40
transitioned to tracheostomy collar | 40
enteral nutrition through jejunostomy feeding tube | 40
left intensive care unit | 40
discharged home | 114
endoscopy surveillance | 114
progression and further extend of disease | 114
bronchoscopies | 1, 8, 17 weeks
tracheoesophageal fistula | 17 weeks
esophageal lumen opening at midway through posterior wall of trachea | 17 weeks
esophagoduodenoscopy | 28 weeks
tracheostomy tube through a combined lumen formed by esophagus and trachea | 28 weeks
double lumen identified with esophagus opening at proximal end of stent | 28 weeks
complete obliteration of stent due to in-growth tissues | 28 weeks
cardiothoracic surgical evaluation | 28 weeks
nutritional optimization | 28 weeks
potential surgical intervention | 28 weeks