84 years old | 0  
    immunocompetent male | 0  
    presented with right inguinal pain | -72  
    presented with fever | -72  
    presented with decreased appetite | -72  
    presented with limited mobility | -72  
    obesity | 0  
    permanent atrial fibrillation | 0  
    apixaban | 0  
    chronic kidney disease stage IIIb | 0  
    distant repaired abdominal aortic aneurysm | 0  
    endovascular graft | 0  
    motor vehicle accident 3 months prior | -2016  
    left knee hemarthrosis | -2016  
    left lower limb cellulitis | -2016  
    cellulitis resolved | -2016  
    hypotensive | 0  
    blood pressure 95/61 mmHg | 0  
    borderline febrile 37.8°C | 0  
    hypoxic | 0  
    oxygen saturation 90% | 0  
    heart rate 75/min | 0  
    weight 114.4 kg | 0  
    alert and oriented | 0  
    cardiovascular examination unremarkable | 0  
    inguinal examination unremarkable | 0  
    ocular examination unremarkable | 0  
    no peripheral stigmata of infective endocarditis | 0  
    cellulitis in left lower limb | 0  
    erythema extending from hemarthrosis scar | 0  
    possible inoculation | 0  
    acute on chronic renal impairment | 0  
    creatinine 111 μmol/L | 0  
    creatinine 149 μmol/L 2 months prior | -1440  
    albumin 32 g/L | 0  
    total bilirubin 18 μmol/L | 0  
    creatinine kinase 72 U/L | 0  
    aspartate aminotransferase 14 U/L | 0  
    alanine transferase 10 U/L | 0  
    white cell count 8.7 × 109/L | 0  
    neutrophil count 7.24 × 109/L | 0  
    lymphocytes 0.66 × 109/L | 0  
    pH 7.45 | 0  
    HCO3 22 mmol/L | 0  
    lactate 2.3 mmol/L | 0  
    coagulation profile unremarkable | 0  
    lymphocyte subsets unremarkable | 0  
    immunoglobulin subsets unremarkable | 0  
    HIV serology unremarkable | 0  
    C-reactive protein 95 mg/L | 0  
    C-reactive protein 150 mg/L | 48  
    SOFA score 3 | 24  
    CT angiography negative for acute aortic syndrome | 0  
    CT angiography negative for vascular graft involvement | 0  
    IV flucloxacillin 2 g | 0  
    IV gentamicin 420 mg | 0  
    IV vancomycin 1 g | 0  
    IV crystalloid fluid resuscitation | 0  
    three liters of fluid resuscitation | 0  
    required metaraminol infusion | 0  
    MAP >65 mmHg | 0  
    metaraminol infusion 0.5 mg/h | 0  
    admitted to intensive care unit | 0  
    intensive care stay 3 days | 72  
    hypoxia improved | 0  
    blood cultures positive for S. schleiferi ssp. coagulans | 24  
    Gram stain identification | 24  
    matrix-assisted laser desorption/ionization time-of-flight mass spectrometry | 24  
    urease-positive | 24  
    coagulase-positive | 24  
    blood cultures repeatedly positive | 24  
    IV piperacillin/tazobactam 4.5 g 6 h | 24  
    IV vancomycin 2 g loading dose | 24  
    IV vancomycin 1 g twice daily | 24  
    antimicrobial susceptibilities returned | 24  
    IV flucloxacillin | 24  
    transthoracic echocardiography unremarkable | 24  
    transesophageal echocardiography unremarkable | 24  
    CT-PET indicated FDG uptake in left iliac graft | 72  
    SUVmax 4.9 | 72  
    history of exposure to pet Maltese terrier's otorrhea | -168  
    canine's otitis externa preceded by a week | -168  
    canine treated with topical miconazole nitrate | -168  
    canine treated with topical prednisolone acetate | -168  
    canine treated with topical polymyxin B | -168  
    canine licked the patient | -168  
    exposure to canine's otorrhea during antimicrobial application | -168  
    left knee hemarthrosis | 0  
    canine aural samples posttreatment positive for Staphylococcus intermedius group | -168  
    vascular surgical opinion obtained | 72  
    multidisciplinary team discussion | 72  
    indefinite antimicrobial suppression with oral flucloxacillin | 72  
    IV flucloxacillin 2 g 4 h for 6 weeks | 72  
    pulmonary edema secondary to fluid resuscitation | 72  
    diuresis with daily furosemide | 72  
    discharged | 72  
    outpatient parental antimicrobial therapy | 72  
    oral antimicrobial suppression | 72