sudden development of fecal incontinence | -12
left hemiplegia | -12
dextroversion | -12
dysarthria | -12
vomiting | -12
transported to the emergency department | -1.33
impaired consciousness | 0
Glasgow coma scale score of 12 | 0
systolic blood pressure, 91 mmHg | 0
respiratory rate, 24/min | 0
oxygen saturation of arterial blood (SpO2), 86% | 0
poor oral hygiene | 0
diminished breath sounds on the left side | 0
coarse crackles in the right lung | 0
decrease in breath sounds in the front of the chest | 0
respiratory condition deteriorated rapidly | 0
endotracheal intubation | 0.67
mechanical ventilation initiated | 0.67
bilateral infiltration on chest CT | 0.67
admitted to the intensive care unit (ICU) | 0.67
leukocyte count (1900/μL) | 0
mildly elevated C-reactive protein (CRP) level (3.6 mg/dL) | 0
respiratory failure with a partial pressure of oxygen in arterial blood (PaO2) of 64 mmHg | 0
hepatorenal function normal | 0
extensive infiltration shadows on chest radiography | 0
hematoma extending from the right basal ganglia and putamen to the thalamus on head CT | 0
consolidations admixture with ground-glass opacities on chest CT | 0
A-DROP score indicated ICU admission | 0
antigen test for coronavirus disease 2019 negative | 0
sputum culture showed Streptococcus agalactiae and Klebsiella oxytoca | 12
management in the ventilator mode started with meropenem and levofloxacin | 12
prednisolone started at 1 mg/kg/day | 12
infiltration shadows improved by Day 12 | 288
extubated on Day 12 | 288
transferred to the Department of Neurosurgery on Day 22 | 528
transferred to a rehabilitation hospital for sequelae of stroke | 528