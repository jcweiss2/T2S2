61 years old | 0
    male | 0
    T-cell lymphoma | -2016
    chemotherapy | -2016
    deep venous thrombosis | -2016
    pulmonary embolism | -2016
    therapeutic anticoagulation | -2016
    typhlitis | -2016
    terminal ileum infiltration | -2016
    cecum infiltration | -2016
    pulmonary involvement | -2016
    bilateral pleural effusions | -2016
    ground-glass opacification | -2016
    alveolar opacities | -2016
    respiratory failure | -2016
    sepsis | -2016
    acute tubular necrosis | -2016
    obtundation | 0
    fever | 0
    chills | 0
    diarrhea | 0
    extensive vasogenic edema in right frontal region | -24
    extensive vasogenic edema in left parietal region | -24
    extensive vasogenic edema in bilateral temporal regions | -24
    extensive vasogenic edema in left cerebellar region | -24
    unresponsive | 0
    agonal breathing | 0
    unequal pupils | 0
    herniation syndrome concern | 0
    neurointensive care unit admission | 0
    noncontrast CT head lesions left temporal | 0
    noncontrast CT head lesions left basal ganglia | 0
    noncontrast CT head lesions left occipital lobe | 0
    noncontrast CT head lesions right temporal lobe | 0
    surrounding vasogenic edema | 0
    lesions in superior cerebellum | 0
    lesions in brainstem | 0
    extensive edema | 0
    multifocal lymphoma suspicion | 0
    differential diagnoses: cerebral toxoplasmosis | 0
    differential diagnoses: neurocysticercosis | 0
    differential diagnoses: multiple abscesses | 0
    no acute hemorrhage | 0
    no midline shift | 0
    contrast-enhanced MRI brain lesions | 0
    contrast-enhanced MRI cervical spine lesions | 0
    contrast-enhanced MRI thoracic spine lesions | 0
    leptomeningeal enhancement thoracic spine | 0
    osseous hyperdensities T6 | 0
    osseous hyperdensities T8 | 0
    osseous hyperdensities T12 | 0
    osseous hyperdensities L1 | 0
    osseous hyperdensities L4 | 0
    osseous hyperdensities L5 | 0
    intradural extramedullary lesion C7-T1 | 0
    right temporal craniotomy | 0
    biopsy under stereotactic navigation | 0
    steroids not administered | 0
    ALK-positive anaplastic large T-cell lymphoma diagnosis | 0
    tumor cells positive for CD4 | 0
    tumor cells positive for CD45 | 0
    tumor cells positive for CD30 | 0
    reactive astrocytosis | 0
    cavitation | 0
    rarefaction of brain parenchyma | 0
    postoperative day 1 unresponsiveness | 24
    postoperative day 1 critical illness | 24
    positive IgG antibody against toxoplasmosis | 24
    sulfadiazine treatment | 24
    pyrimethamine treatment | 24
    postoperative day 3 pupils 2mm | 72
    postoperative day 3 nonreactive pupils | 72
    communicating hydrocephalus | 72
    external ventricular catheter placement | 72
    ICP monitoring | 72
    therapeutic ventricular drainage | 72
    head of bed elevation | 72
    blood pressure control | 72
    deep sedation | 72
    elevated ICPs | 72
    postoperative day 7 loss of brainstem reflexes | 168
    bilateral fixed pupils | 168
    bilateral dilated pupils | 168
    severe thrombocytopenia | 168
    multiple platelet transfusions | 168
    hemodynamic instability | 168
    norepinephrine support | 168
    phenylephrine support | 168
    epinephrine support | 168
    vasopressin support | 168
    care withdrawal | 168
    patient expired | 168

<|eot_id|>