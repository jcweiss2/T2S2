68 years old | 0
male | 0
admitted to the hospital | 0
tachypnea | -720
increased FIO2 requirements | -720
endotracheal intubation | -720
mechanical ventilation | -720
morbid obesity | 0
systemic arterial hypertension | 0
diabetes mellitus | 0
chronic lung disease | 0
heavy smoking history | 0
ramipril | 0
amlodipine | 0
metformin | 0
metoprolol | 0
no recent corticosteroids therapy | 0
no immunosuppressive agents | 0
blood pressure 86/52 mm Hg | 0
heart rate 104 beats/min | 0
respiratory rate 24 breaths/min | 0
temperature 37 °C | 0
bilateral rales | 0
wheezing | 0
WBC count 16.4 × 10^3/mm^3 | 0
ALT level 119 U/L | 0
LDH level 488 U/L | 0
BUN level 36 mg/DL | 0
creatinine level normal | 0
cardiac enzymes normal | 0
coagulation profile normal | 0
HIV test negative | 0
arterial blood gas | 0
pH 7.24 | 0
pCO2 level 69 mm Hg | 0
PaO2 level 67 mm Hg | 0
chest X-ray | 0
bilateral increased interstitial markings | 0
left retrocardiac consolidation | 0
chest CT | 0
bilateral ground-glass opacities | 0
no pulmonary embolism | 0
venous Doppler ultrasound | 0
no deep venous thrombosis | 0
electrocardiogram | 0
sinus tachycardia | 0
no ST-segment or T-wave abnormalities | 0
transthoracic echocardiogram | 0
normal left ventricular ejection fraction | 0
normal right ventricular systolic function | 0
no pulmonary hypertension | 0
empiric intravenous antimicrobial therapy | 0
vancomycin | 0
cefepime | 0
azithromycin | 0
vasopressors | 0
norepinephrine | 0
septic shock | 0
community-acquired pneumonia | 0
blood cultures negative | 0
respiratory cultures negative | 0
Legionella urinary antigens negative | 0
Streptococcus pneumoniae urinary antigens negative | 0
serum cryptococcal antigen negative | 0
procalcitonin level 0.25 ng/mL | 0
(1-3)-β-D-glucan assay 32 pg/mL | 0
ICU clinical course complicated | 0
persistently increased FIO2/PEEP requirements | 0
ARDS | 0
decreased PaO2/FIO2 ratio | 0
worsening bilateral infiltrates | 0
increased vasopressors requirements | 0
acute kidney injury | 0
optimal sedation | 0
fentanyl | 0
propofol | 0
neuromuscular blocking agent | 0
cisatracurium | 0
epoprostenol | 0
refractory hypoxemia | 0
extracorporeal membrane oxygenation | 0
inappropriate | 0
plateau pressures < 35 cm H2O | 0
BAL result positive for Pneumocystis jirovecii | 144
CMV antigenemia negative | 144
all serum immunoglobulin levels normal | 144
complement component 3 diminished | 144
complement component 4 diminished | 144
CH50 levels diminished | 144
repeated HIV test non-reactive | 144
T-lymphocytes cell count 97 cells/µL | 144
absolute lymphocytes cell count 377 × 10^3/µL | 144
intravenous antimicrobial therapy | 144
trimethoprim-sulfamethoxazole | 144
steroids | 144
methylprednisone | 144
repeated chest CT | 168
diffuse ground-glass opacities | 168
severe pneumomediastinum | 168
pneumopericardium | 168
bilateral pneumothorax | 168
patient’s clinical condition worsened | 168
withdrawal of artificial life support | 336
patient expired | 336