67 years old | 0
male | 0
diabetes | 0
hypertension | 0
dyslipidemia | 0
left foot pain | -48
left foot swelling | -48
ulcer in the plantar aspect | -48
pus discharge | -48
fever | -48
generalized weakness | -48
admitted to the hospital | 0
febrile | 0
tachycardic | 0
left foot swelling | 0
hotness | 0
redness | 0
tenderness | 0
left plantar ulcer | 0
pus discharge | 0
necrotic base | 0
folly catheter inserted | 0
pus in urine | 0
WBC 15.5 | 0
hemoglobin 7.9 | 0
CRP 41 | 0
potassium 5.5 | 0
sodium 130 | 0
random blood glucose 327 | 0
urine showed numerous WBC and RBC | 0
left plantar ulcer debridement | 0
daily dressing | 0
intravenous antibiotic | 0
sudden onset severe abdominal pain | 72
abdominal pain in suprapubic region | 72
fever | 72
vomiting | 72
abdomen distended | 72
abdomen tense | 72
abdomen tender | 72
abdominal CT scan | 72
moderate pneumoperitoneum | 72
moderate abdomino-pelvic free fluid | 72
hollow viscus perforation | 72
diffuse haziness in the mesentery | 72
moderate dilatation of the small bowel loops | 72
Foley’s catheter balloon seen in situ | 72
partially distended urinary bladder | 72
perforated viscus | 72
exploratory laparotomy | 96
moderate intra-abdominal turbid fluid collection | 96
pockets of pus in the pelvis | 96
pockets of pus in the right paracolic gutter | 96
dilated congested bowel loop | 96
edema of the mesentery | 96
urinary bladder perforation | 96
inflamed mucosa | 96
pus coming from inside the urinary bladder | 96
lavage of the peritoneal cavity | 96
biopsies taken from the edges of the perforation | 96
refreshed edges of the perforation | 96
water tight repair | 96
suprapubic catheter inserted | 96
Foley’s catheter inserted | 96
nonspecific inflammation of bladder wall | 120
no evidence of malignancy | 120
post-operative recovery | 120
transferred to the surgical ward | 168
started oral fluids | 168
full diet commenced | 240
intravenous antibiotics continued | 240
discharged from the hospital | 240