65 years old | 0
male | 0
autoimmune hepatitis | 0
hypertension | 0
hyperlipidemia | 0
benign prostatic hypertrophy | 0
admitted to ICU | 0
severe symptomatic hypotonic hyponatremia | 0
furosemide | 0
allopurinol | 0
prazosin | 0
folic acid | 0
ursodiol | 0
pantoprazole | 0
prednisolone | 0
DLBCL of liver | -720
cyclophosphamide | 0
rituximab | 0
dexamethasone | 0
tumor lysis syndrome | 0
renal failure | 0
hemodialysis | 0
volume overload | 0
respiratory failure | 0
intubation | 0
mechanical ventilation | 0
extubated | 0
transferred to oncology service | 0
chest CT | 432
PEA arrest | 432
central airway obstruction | 432
blood clots | 432
emergent intubation | 432
return of spontaneous circulation | 435
cachectic | 432
fever | 432
temperature 38.2°C | 432
pulse 72/min | 432
blood pressure 107/61 mmHg | 432
respiratory rate 21 | 432
oxygen saturation 97% | 432
FiO2 50% | 432
dried blood in oropharynx | 432
bloody secretions | 432
anasarca | 432
WBC 3.8 10^3/uL | 432
hemoglobin 9.5 g/dL | 432
BUN 56 mg/dL | 432
creatinine 1.69 mg/dL | 432
thick-walled cavitary lesion | 408
air fluid level | 432
bronchoscopy | 432
extensive blood clots | 432
thick mucus | 432
CT pulmonary angiography | 432
saccular contrast-enhancing lesion | 432
PAP | 432
PM | 432
Mucor | 432
isavuconazonium | 432
embolization | 480
no further hemoptysis | 480
irreversible anoxic brain injury | 480
nonresponsive | 480
renal failure worsened | 480
forgo hemodialysis | 480
forgo cardiopulmonary resuscitation | 480
passed away | 744