31 years old | 0 | 0 
female | 0 | 0 
SLE | -8760 | 0 
lupus nephritis | -8760 | 0 
prior stroke | -8760 | 0 
intravenous drug use | -8760 | 0 
cardiogenic shock | 0 | 0 
mental status changes | 0 | 0 
elevated jugular venous pressure | 0 | 0 
prominent v wave | 0 | 0 
body temperature 36.3°C | 0 | 0 
blood pressure 95/66 mm Hg | 0 | 0 
heart rate 94 beats/min | 0 | 0 
hemoglobin 10.3 g/dL | 0 | 0 
white blood cell count 18.9 × 10^9/L | 0 | 0 
platelet count 64 × 10^9/L | 0 | 0 
international normalized ratio 3.6 | 0 | 0 
creatinine level 1.7 mg/dL | 0 | 0 
drug studies positive for narcotics | 0 | 0 
drug studies positive for cannabis | 0 | 0 
antiphospholipid serology normal | 0 | 0 
blood cultures negative | 0 | 0 
intravenous antibiotics | 0 | 24 
broad-spectrum intravenous antibiotics | 0 | 24 
NBTE | -168 | 0 
mitral valve replacements | -168 | -168 
aggressive immunosuppression | -168 | -168 
anticoagulation | -168 | -168 
mitral valve prosthesis dehiscence | 0 | 0 
severe perivalvular regurgitation | 0 | 0 
annular pseudoaneurysm | 0 | 0 
left atrial thrombus | 120 | 120 
surgical clot removal | 120 | 120 
recurrent left atrial thrombus | 120 | 168 
extracorporeal membrane oxygenation | 24 | 168 
multiple blood product transfusions | 24 | 168 
left ventricular ejection fraction 25% | 24 | 168 
sluggish flow in the left atrium | 24 | 168 
death | 168 | 168 
autopsy declined | 168 | 168 
transthoracic echocardiography | 0 | 0 
transesophageal echocardiography | 0 | 0 
three-dimensional imaging | 0 | 0 
color Doppler | 0 | 0 
valvular surgery | 0 | 168 
valvular reconstruction | 24 | 168 
mitral valve annulus reconstruction | 24 | 168 
bioprosthesis | 24 | 168 
bovine pericardium | 24 | 168 
left atrial dome reconstruction | 24 | 168 
interatrial septal incision reconstruction | 24 | 168 
postoperative TEE | 24 | 168 
layered thrombus in the left atrium | 120 | 120 
thrombus reaccumulation | 120 | 168 
extracorporeal membrane oxygenation withdrawal | 168 | 168