41 years old | 0
male | 0
morbid obesity | 0
admitted to the hospital | 0
painful bilateral oedema of lower legs | 0
generalized abdominal pain | 0
liver cirrhosis | -672
excessive alcohol abuse | -672
hepatitis C infection | -672
portal hypertension | -672
oesophageal varices | -672
febrile | 0
bilateral pitting oedema | 0
superficial pre-tibial abrasions | 0
capillary refill time normal | 0
distal pulses present | 0
abdominal examination unremarkable | 0
respiratory examination unremarkable | 0
cardiovascular examination unremarkable | 0
neurological examination unremarkable | 0
low haemoglobin | 0
platelet count low | 0
albumin low | 0
bilirubin elevated | 0
CRP elevated | 0
INR elevated | 0
lactate elevated | 0
liver enzymes normal | 0
Child's B case of cirrhosis | 0
blood cultures performed | 0
swab of left leg performed | 0
treatment started with flucloxacillin and benzylpenicillin | 0
left leg swelling increased | 24
overlying skin erythematous | 24
tender to touch | 24
induration | 24
blistering | 24
CRP increased | 24
ciprofloxacin and cephazolin started | 24
left leg duplex ultrasound performed | 24
severe oedema below knee | 24
large knee joint effusion | 24
no deep vein thrombosis | 24
CT scan of legs performed | 24
bilateral knee joint effusions | 24
non-specific synovitis | 24
no necrotizing fasciitis | 24
A. baumannii isolated from blood cultures | 48
A. baumannii resistant to amoxicillin, amoxicillin/clavulanate, ceftriaxone, and ceftazidime | 48
A. baumannii sensitive to co-trimoxazole, gentamycin, meropenem, ciprofloxacin, and ticarcillin/clavulanate | 48
antibiotic regime changed to meropenem and vancomycin | 48
conservative management of lower limbs continued | 48
referred to reconstructive and orthopaedic surgeons | 48
MRI scan of lower legs performed | 72
extensive subcutaneous oedema | 72
mild to moderate subcutaneous oedema | 72
moderate bilateral joint effusions | 72
cellulitic changes | 72
extensive myositis | 72
possible fasciitis | 72
lincomycin added to therapy | 72
fever | 96
left leg surgically explored | 96
no evidence of necrotizing fasciitis | 96
no evidence of compartment syndrome | 96
extensive subcutaneous oedema | 96
circumferential debridement of fat necrosis and muscle | 96
washout of left leg wound | 96
VAC dressing applied | 96
antibiotics continued | 96
ventilated post-operatively | 96
noradrenaline infusion started | 96
cultures from left leg subcutaneous tissue confirmed A. baumannii | 96
antibiotic regime changed to ciprofloxacin, meropenem, and lincomycin | 96
vancomycin ceased | 96
further surgical debridement performed | 144
necrotic circumferential subcutaneous fat | 144
circumferential debridement of subcutaneous tissue | 144
washout with hydrogen peroxide | 144
new VAC dressing applied | 144
histopathology revealed epidermal and dermal infarction | 144
focal fat necrosis | 144
acute inflammation | 144
no histological evidence of fasciitis | 144
antibiotic management tailored to meropenem and ciprofloxacin | 144
further surgical procedures performed | 192
VAC dressing changed | 192
wound reviewed | 192
necrosis along wound edges | 192
minor debridement performed | 192
VAC dressing replaced | 192
wound reviewed | 240
significant improvement | 240
small areas of necrotic tissue | 240
minor debridement performed | 240
samples sent for microscopy and culture | 240
wound washed with hydrogen peroxide | 240
clinically jaundiced | 240
worsening hepatic and renal function | 240
condition deteriorated | 240
hepatic failure | 240
circulatory failure | 240
respiratory failure | 240
haematological failure | 240
blood glucose levels fluctuated | 240
inotrope dependent | 240
insulin required | 240
decision to palliate made | 336
died | 336