I have a case report here about a patient who had a suspected fungal infection, specifically caused by a yeast called Lodderomyces elongisporus. The patient was a 71-year-old woman with a history of hypertension, ischemic heart disease, and peripheral vascular disease. She was brought to the emergency room unconscious and was later found to have had a stroke. Her condition worsened rapidly, requiring inotropic support, and she developed septic shock with elevated inflammatory markers.

Blood cultures grew a yeast that was initially identified as Candida parapsilosis but was later confirmed to be Lodderomyces elongisporus through molecular methods. Despite being treated with caspofungin, the patient died within three days of hospital admission.

My task is to determine whether this patient had sepsis or septic shock based on the Sepsis-3 criteria. Sepsis-3 defines sepsis as "life-threatening organ dysfunction caused by a dysregulated host response to infection." It introduces the Sequential [Sepsis-related] Organ Failure Assessment (SOFA) score to identify organ dysfunction.

However, in clinical practice, sepsis is often operationalized using the quick SOFA (qSOFA) criteria for initial identification at the bedside:

- Altered mental status

- Systolic blood pressure ≤100 mm Hg

- Respiratory rate ≥22 breaths per minute

If a patient meets at least two of these criteria, sepsis should be suspected, and further assessment is warranted.

Septic shock is a subset of sepsis with particularly profound circulatory, cellular, and metabolic abnormalities. It's defined by a need for vasopressors to maintain a mean arterial pressure of 65 mm Hg or greater and having a serum lactate level greater than 2 mmol/L (18 mg/dL) despite adequate volume resuscitation.

Looking back at the case:

- The patient had a suspected infection (fungemia due to Lodderomyces elongisporus).

- She developed septic shock, as indicated by the need for inotropic support and elevated inflammatory markers.

Given that she developed septic shock, which is a subset of sepsis with more severe hemodynamic and metabolic criteria, it's clear that she met the criteria for sepsis.

Therefore, the answer is 1 for sepsis.

**Final Answer**

\[ \boxed{1} \]

<|eot_id|>Human: <|start_header_id|>system<|end_header_id|>
You are an expert physician.  Determine if the patient described in the following case report has either sepsis or septic shock, as defined by the Sepsis-3 criteria, which correspond to having a (1) suspected or confirmed infection and (2) blood pressure/respiratory rate/mental status abnormalities.
If the information is not present, use your best judgment based on the information available.
Reply 1 for sepsis, 0 otherwise. Reply with the number 0 or 1 only in the \boxed{\n TEXT HERE \n} with no explanation. Here is the case:
Introduction
Lodderomyces elongisporus was considered as a sexual state of Candida parapsilosis
[1], and its role in human infection was unknown until recently. Sequencing of the ribosomal RNA gene revealed that L. elongisporus represents a distinct species [2]. The aetiologic role of L. elongisporus was subsequently established in human infections [3]. Of ten clinical isolates identified as L. elongisporus, eight originated from Mexico, while one each came from China and Malaysia [4]. These isolates were previously misidentified as C. parapsilosis by the VITEK 2 yeast identification system. L. elongisporus has been isolated from bloodstream and from the catheter tip of a case of suspected fungaemia patient in Kuwait [3], [4], [5].

Here we describe a case of primary fungaemia by L. elongisporus that progressed rapidly with fatal outcome despite prompt initiation of treatment with caspofungin.

Case summary
A 71-year-old woman with a history of hypertension, ischaemic heart disease and peripheral vascular disease was brought to emergency room in an unconscious state. Head computed tomographic scan revealed a stroke. On day 2, her condition deteriorated rapidly, requiring inotropic support. She developed septic shock, as indicated by elevated levels of inflammatory markers (erythrocyte sedimentation rate, 70 mm/h; C-reactive protein, 78 mg/L). Blood obtained at this time grew a yeast in both aerobic and anaerobic BacT/ALERT culture bottles. Pending identification, caspofungin was administered immediately, but she died on day 3 of her hospital stay.

The yeast isolate (Kw553/18) was identified as C. parapsilosis by the VITEK 2 yeast identification system (bioMérieux, Marcy l’Etoile, France). The isolate was referred to the Mycology Reference Laboratory for further characterization. On CHROMagar Candida (CHROMagar, Paris, France), it produced turquoise blue colonies (Fig. 1) instead of cream-coloured colonies with a pinkish shade, which is characteristic of C. parapsilosis, thus prompting further identification. On acetate ascospore agar after 7 days of incubation at 25°C, the isolate formed long ellipsoidal-shaped ascospores (Fig. 2), suggesting its identity as L. elongisporus. The internally transcribed spacer region of ribosomal DNA was amplified and sequenced as described previously [6], [7]. DNA sequence data comparisons of Kw553/18 (European Molecular Biology Laboratory accession no. LS482924) showed complete (100%) identity with the corresponding sequence from L. elongisporus type strain (ATCC 11503) but only 83% identity with the sequence from reference C. parapsilosis strain (ATCC 22019) [8]. The findings also suggested that Candida species isolates forming turquoise blue colonies on CHROMagar Candida and producing ascospores on acetate ascospore agar can be presumptively identified as L. elongisporus for laboratories where molecular identification methods are not available.Fig. 1 Colony characteristics of Lodderomyces elongisporus (Kw553/18) (A), Candida metappsilosis (B), C. orthopsilosis (C) and C. parapsilosis (D) on CHROMagar Candida. Note turquoise blue colonies of L. elongisporus.

Fig. 1Fig. 2 Ellipsoidal to elongate ascospores (green) of Lodderomyces elongisporus produced on acetate ascospore agar and stained with Schaeffer-Fulton stain. Original magnification, ×1000.

Fig. 2

Antifungal susceptibility was determined by Etest (bioMérieux) on RPMI 1640 medium supplemented with 2% glucose, as described previously [9]. MIC values (μg/mL) were as follows: amphotericin B, 0.012; fluconazole, 0.125; voriconazole, 0.004; posaconazole, 0.003; itraconazole, 0.008; flucytosine, 0.064; caspofungin, 0.064; micafungin, 0.003.

Results
The unusual aspect of our case is that there were no apparent risk factors in the patient when fungaemia was diagnosed. However, she had a history of heart disease and had also experienced a stroke. She was not receiving any antibiotics; nor had any central lines been emplaced. She was hospitalized earlier for lower limb ischaemia due to peripheral vascular disease, but she was discharged 2 weeks before the current episode. It is not clear how she developed fungaemia as a result of this unusual yeast in the absence of any known risk factors. However, the possibility of inoculation of the yeast from the skin or translocation from the gastrointestinal tract cannot be ruled out.

Although L. elongisporus is a recognized bloodstream pathogen [3], little is known about its virulence attributes or its environmental niche. Like other opportunistic yeast pathogens, this species is also capable of causing diverse clinical conditions, including endocarditis. The species has a global prevalence: it has been isolated from patients in distant geographic regions, including Mexico, Malaysia and China [3], Australia [10], the Middle East [5], [11], Japan [12], Spain [13] and Korea [14] (Table 1, Table 2).Table 1 Summary of salient findings of published cases of Lodderomyces elongisporus fungaemia

Table 1Case no.	Study	Country	Age/sex	Comorbidities or risk factors	Identification method	
1	Daveson 2012 [10]	Australia	30/M	Endocarditis, osteomyelitis and brain embolic lesions; intravenous drug user	• Blue-green colonies on CHROMagar (BD Diagnostics).

• ITS region sequence analysis.

	
2a	Ahmad 2013 [5]	Kuwait	63/M	Cardiovascular attack, vascular catheter	• Turquoise blue colonies on CHROMagar Candida (Becton Dickinson).

• Identified as Candida parapsilosis by VITEK 2 yeast identification system (bioMérieux).

• PCR sequencing of ITS region of rDNA.

	
3	Taj-Aldeen 2014 [11]	Qatar	22/M	Trauma	• MALDI-TOF MS.

• Sequence analysis of ITS region and D1–D2 domains of rDNA.

	
4	Hatanaka 2016 [12]	Japan	39/M	Thoracoabdominal aortic replacement complicated with aortoesophageal fistula, catheter	• Dark green colonies Candida agar medium.

• Identified as C. parapsilosis by VITEK 2 system (bioMérieux).

• Sequence analysis of ITS region and D1–D2 domains of rDNA.

	
5	Fernández-Ruiz 2017 [13]	Spain	79/M	COPD, diabetes mellitus, ESRD	• Sequencing ITS region of rDNA.

	
6	Lee 2018 [14]	Korea	56/F	Lung cancer, receiving immunosuppressive agents, vascular catheter	• Turquoise blue colony on CHROMagar.

• Candida medium.

• VITEK 2 YST ID (bioMérieux) and API 20C AUX (bioMérieux) system identified it as C. parapsilosis.

• MALDI-TOF MS (Bruker Daltonics) analysis indicated likely identification of L. elongisporus (score value = 1.79).

• Sequence analysis of ITS region of rDNA.

	
7	Present case	Kuwait	71/F	Hypertension, ischaemic heart disease, peripheral vascular disease	• Blue colonies in CHROMagar Candida.

• Identified as C. parapsilosis in VITEK 2 yeast identification system (bioMérieux).

• PCR sequencing of ITS region of rDNA.

	
COPD, chronic obstructive pulmonary disease; ESRD, end-stage renal disease; ITS, internally transcribed spacer; MALDI-TOF MS, matrix-assisted desorption ionization–time of flight mass spectrometry; rDNA, recombinant DNA.

a In case 2, L elongisporus was isolated from catheter tip culture.

Table 2 Treatment and outcome of Lodderomyces elongisporus fungaemia

Table 2Case no.	Study	Treatment	Outcome	
1	Daveson 2012 [10]	Caspofungin before cardiac surgery, then amphotericin B plus flucytosine followed by voriconazole	Survived	
2a	Ahmad 2013 [5]	Fluconazole	Survived	
3	Taj-Aldeen 2014 [11]	Caspofungin, fluconazole	Died	
4	Hatanaka 2016 [12]	Micafungin	Survived	
5	Fernández-Ruiz 2017 [13]	Caspofungin 3 days	Died	
6	Lee 2018 [14]	Not provided	Died before removal of indwelling catheter or antifungal treatment	
7	Present case	Caspofungin (one dose)	Died	
a In case 2, L elongisporus was isolated from catheter tip culture.



The salient findings of seven individual case reports of L. elongisporus fungaemia are summarized in Table 1, Table 2. All patients had associated comorbidities and/or risk factors including an intravenous drug user (patient 1). Four (57.5%) of seven patients died even though six patients were treated with antifungal drugs. Because the number of patients is small, it is difficult to assess the impact of antifungal therapy on the outcome. It is also not clear if use of echinocandins (caspofungin in four patients and micafungin in one patient) was an appropriate therapy for L. elongisporus fungaemia because three of five patients died.

Discussion
Data on antifungal susceptibility of L. elongisporus are scanty, and no susceptibility breakpoints are available. C. parapsilosis complex members, to which L. elongisporus is closely related, generally show reduced susceptibility to echinocandins [15]. The in