67 years old | 0
female | 0
admitted to the hospital | 0
fever | -96
chills | -96
cough | -96
dyspnea | -96
diabetes mellitus | 0
temperature of 38.9°C | 0
mild icterus | 0
bilateral rhonchi | 0
crepitations on lung auscultation | 0
no tenderness over right hypochondrial region | 0
raised white blood cell count (10,400/mL) | 0
90.2% neutrophils | 0
hemoglobin level of 11.0 g/dL |1 0
platelet count of 81,000/μL | 0
aspartate aminotransferase level of 86 units/L | 0
alanine aminotransferase of 78 units/L | 0
high total bilirubin (49.3 μmol/L) | 0
high blood glucose (18.4 mmol/L) | 0
acute kidney injury | 0
blood urea nitrogen 24 mg/dL | 0
creatinine of 1.7 mg/dL | 0
chest CT scan showing SPE | 0
multiple peripheral nodules in both lungs | 0
wedge-shaped peripheral infiltrative lesions abutting pleura | 0
bilateral pleural effusions | 0
liver mass | 0
transthoracic echocardiography showing mild tricuspid regurgitation | 0
no vegetations on heart valves | 0
intravenous imipenem | 0
fever worsened | 0
chills worsened | 0
dyspnea worsened | 0
contrast-enhanced abdominal CT | 48
large liver abscess without gas formation | 48
pneumocardia with air within right ventricle | 48
supine Trendelenburg position | 48
100% oxygen administered | 48
admission to telemetry unit | 48
liver abscess drained | 48
continued intravenous imipenem | 48
symptoms improved gradually | 72
transthoracic echocardiography no air in heart | 72
positive blood cultures | 72
positive pus culture from liver abscess | 72
Klebsiella pneumoniae | 72
discharged | 600
follow-up at 10 months | 7200
