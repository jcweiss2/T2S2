62 years old | 0
male | 0
admitted to the hospital | 0
fever | -48
high-grade fever | -48
arthralgia | -48
generalized malaise | -48
hypotension | -48
shock | -48
systolic blood pressure 72 mmHg | -48
heart rate 110 beats per minute | -48
pain in the lateral aspect of the right elbow | -48
tachypneic | 0
not in shock | 0
BP 102/66 mmHg | 0
HR 114 beats per minute | 0
respiratory rate 28 breaths per minute | 0
febrile 38.5°C | 0
required oxygen | 0
oxygen saturation 94% on 3 L/min cannula | 0
erythematous and visibly swollen right elbow | 0
tenderness on palpation | 0
entered a state of shock | 0
disseminated intravascular coagulation | 0
multiple organ failure | 0
intensive care | 0
Streptococcus pyogenes in blood cultures | 0
fasciotomy and debridement for necrotizing fasciitis | 0
STSS diagnosed | 0
intubation | 0
vasopressors | 0
antibiotics | 0
fluid management | 0
ventilation support | 0
afebrile on day 15 | 360
high-grade fever on day 34 | 816
hypotension on day 34 | 816
tachycardia on day 34 | 816
leukocytosis on day 34 | 816
evidence of MOF on day 34 | 816
vasopressors on day 34 | 816
abdominal CT demonstrated left IPA | 816
Klebsiella pneumoniae in blood cultures | 816
intravenous antibiotics against Klebsiella pneumoniae | 816
MOF improved without drainage | 816
CT-guided drainage of the abscess on day 53 | 1272
culture of the drainage specimen did not grow any bacteria | 1272
drainage tube removed 2 weeks after the procedure | 1596
follow-up abdominal CT confirmed significant shrinkage of the IPA | 1596
rehabilitation | 1596
discharged on foot | 1596
follow-up for more than 2 years | 4320
excellent results in activities of daily living | 4320