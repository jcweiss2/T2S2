33 years old | 0
male | 0
183 cm | 0
94 kg | 0
admitted to the hospital | 0
severe abdominal pain | 0
vomiting | -24
abdominal pain developed | -24
visited another hospital | -24
minor mental deterioration | -24
transferred to the ER | 0
blood pressure 105/63 mmHg | 0
heart rate 69 beats/min | 0
peripheral oxygen saturation 99% | 0
respiratory rate 20 rates/min | 0
body temperature 36.9℃ | 0
arterial blood gas analysis | 0
pH 7.64 | 0
arterial CO2 partial pressure 25.8 mmHg | 0
arterial O2 partial pressure 111.1 mmHg | 0
base excess 8.3 mmol/L | 0
chest radiograph | 0
chest and abdominal CT | 0
blood pressure 83/66 mmHg | 0
heart rate 116 beats/min | 0
intravenous administration of 100 ml of crystalloid fluids | 0
blood pressure 124/88 mmHg | 0
severe increase in stomach volume | 0
stricture in the gastric pylorus and duodenum | 0
unsuccessful insertion of a nasogastric tube | 0
pneumomediastinum | 0
esophageal rupture | 0
right internal jugular vein catheterization | 0
blood pressure 84/44 mmHg | 0
heart rate 113 beats/min | 0
intravenous administration of 300 ml of crystalloid solution | 0
oxygen administration | 0
SpO2 97% | 0
moved to the operating room | 24
fasting time 12 hours | 24
preoperative blood tests | 24
blood urea nitrogen 32 mg/dl | 24
creatinine 2.2 mg/dl | 24
white blood cell 12,400/mm3 | 24
clear consciousness | 24
blood pressure 80/50 mmHg | 24
heart rate 125 beats/min | 24
SpO2 94% | 24
preoxygenation | 24
general anesthesia | 24
endotracheal intubation | 24
mechanical ventilation | 24
pressure control ventilation | 24
desflurane | 24
dopamine | 24
single right lung ventilation | 24
pneumomediastinum | 24
esophageal rupture | 24
desaturation | 24
manual ventilation | 24
SpO2 80% | 24
two-lung ventilation | 24
SpO2 70% | 24
cardiopulmonary resuscitation | 24
epinephrine | 24
bilateral tension pneumothorax | 24
angiocatheter insertion | 24
air leakage | 24
foul smelling brown liquid | 24
SpO2 90% | 24
heart rate 70-80 beats/min | 24
systolic blood pressure 100-120 mmHg | 24
SpO2 94-95% | 24
emergency chest radiograph | 24
chest tube insertion | 24
breath sounds recovery | 24
SpO2 100% | 24
stomach contents gushing out | 24
lung parenchymal damage | 24
left-lung ventilation | 24
right thoracotomy | 24
stomach contents suctioned out | 24
lung irrigation | 24
chemical burn | 24
esophagectomy | 24
esophagogastrostomy | 24
feeding jejunostomy | 24
fluids administration | 24
blood loss | 24
urine output | 24
arterial blood gas analysis | 24
pH 7.429 | 24
arterial CO2 partial pressure 31.3 mmHg | 24
arterial O2 partial pressure 367.7 mmHg | 24
base excess -2.2 mmol/L | 24
single-lumen tube | 24
intensive care unit | 24
mechanical ventilation | 24
fentanyl | 24
sedation | 24
pain control | 24
arterial blood gas analysis | 26
pH 7.43 | 26
arterial CO2 partial pressure 31 mmHg | 26
arterial O2 partial pressure 211 mmHg | 26
base excess -2 mmol/L | 26
SpO2 99% | 26
mechanical ventilation | 48
FIO2 0.4 | 48
arterial blood gas analysis | 48
pH 7.39 | 48
arterial CO2 partial pressure 35 mmHg | 48
arterial O2 partial pressure 169 mmHg | 48
base excess -2.0 mmol/L | 48
SpO2 99% | 48
T-piece | 120
FIO2 0.35-0.50 | 120
extubation | 168
SpO2 97% | 168
oxygen administration | 168
left-side chest tube removal | 264
right-side chest tube removal | 600
discharge | 768