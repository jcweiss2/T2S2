48 years old | 0
male | 0
admitted to the hospital | 0
smoking | -8760
bowel resection | -720
intense headache | -48
abdominal pain | -48
dyspnoea | -168
generalized oedema | -168
asthenia | -168
decrease in urinary output | -168
non-specific abdominal pain | -720
hypotension | -720
elevated plasma lactate levels | -720
haemoconcentration | -720
metabolic acidosis | -720
normal plasma creatine phosphokinase levels | -720
abdominal CT arteriography | -720
intensive haemodynamic support | -720
monitoring | -720
emergent abdominal exploration | -720
bowel resection | -720
diagnosis of non-occlusive mesenteric ischaemia | -720
catheter-related superior vena cava thrombosis | -720
implantation of a vascular access system | -720
parenteral nutrition | -720
hypocoagulation | -720
oliguric acute renal injury | -1092
hypovolaemic shock | -1092
metabolic acidaemia | -1092
intensive care unit admission | -1092
ionotropic support | -1092
renal replacement treatment | -1092
broad spectrum empiric antibiotics | -1092
prodrome of intense headache | -48
prodrome of diffuse abdominal discomfort | -48
physical exercise | -48
heat exposure | -48
haemodynamically unstable | 0
hypotension | 0
heart rate of 120 bpm | 0
generalized oedema | 0
no skin flushing | 0
no urticaria | 0
no focal angioedema | 0
no stridor | 0
no lymphadenopathy | 0
severe metabolic acidaemia | 0
haemoconcentration | 0
elevated Hgb | 0
elevated haematocrit | 0
leucocytosis | 0
uraemia | 0
elevated creatinine | 0
hypoalbuminaemia | 0
elevated BNP | 0
normal troponin level | 0
normal electrocardiogram | 0
normal thoracic x-ray | 0
normal urinary study | 0
normal contrast-enhanced thoracoabdominal CT scan | 0
normal abdominal and renal ultrasound | 0
intensive fluid replacement therapy | 0
haemodynamic stabilization | 0
renal function recovery | 0
inflammatory studies | 0
complete infectious study | 0
diagnosis of idiopathic systemic capillary leak syndrome | 0
prodromes of intense headache | 0
prodromes of abdominal pain | 0
association with previous heat exposure | 0
thyroid function tests | 0
gonadal function tests | 0
adrenal steroid function tests | 0
immune function tests | 0
metabolic function tests | 0
complement studies | 0
C1 esterase inhibitor levels | 0
C1 esterase inhibitor function | 0
cardiac study | 0
transthoracic echocardiography | 0
cardiovascular MRI | 0
whole endoscopic study | 0
monoclonal gamma/lambda gammopathy | 0
immunofixation | 0
serum free light chain assay | 0
bone marrow biopsy | 0
intravenous immunoglobulin | 0
nutritional supplementation | 720
discharged | 720
oedema of the extremities | 1440
fatigue | 1440
partial leaks | 1440
prophylactic treatment with terbutaline | 1440
prophylactic treatment with theophylline | 1440
periodic plasma level evaluations | 1440
avoided physical exercise | 1440
avoided heat exposure | 1440
hospital admissions for acute exacerbation | 2880
subtherapeutic theophylline levels | 2880
prophylactic administration of IVIG | 2880
good results | 4320