60 years old | 0
male | 0
presented to King Khalid University Hospital | 0
erythroderma | -12960
erythematous lesions | -43440
pruritus | -43440
oral prednisolone | -43440
oral cyclosporine | -43440
confluent lichenified erythromelanotic plaques | 0
thick plate of greasy scales | 0
no lymph node enlargement | 0
bilateral lower lid ectropion | 0
skin punch biopsies taken | 0
epidermotropism of atypical lymphocytes | 0
lymphocytic band infiltrate | 0
dermal fibrosis | 0
negative immunofluorescence study | 0
CD3 positive | 0
CD45RO positive | 0
CD4 negative | 0
CD8 negative | 0
CD7 negative | 0
CD30 positive | 0
normal peripheral blood count | 0
no Sézary cells | 0
flow cytometry negative | 0
CT scan abdomen pelvis | 0
enlarged lymph nodes | 0
CT scan chest | 0
no lymphadenopathy | 0
lymph node biopsy | 0
large atypical cells | 0
negative clonal T-cell rearrangement | 0
diagnosis of double-negative CD4/CD8 MF | 0
referred to hematology oncology unit | 0
septic shock | 288
admitted to intensive care unit | 288
passed away | 360
misdiagnosed as severe eczema | -43440
erythema gyratum repens-like MF | 0
purpuric MF | 0
ichthyosiform MF | 0
complete response to psoralen plus UVA | 0
partial response to phototherapy | 0
indolent course | 0
aggressive behavior | 0
large cell transformation | 0
metastasis | 0
responded partially to treatment | 0
died 5 years after symptoms | 0
died 45 days after diagnosis | 0
