20 years old | 0
male | 0
admitted to the hospital | 0
abdominal pain | -144
watery diarrhoea | -144
nausea | -144
vomiting | -144
fever | -144
chills | -144
cough | -144
shortness of breath | -144
colitis | -144
prescribed oral ciprofloxacin | -144
prescribed metronidazole | -144
achy pain | -144
diffuse pain | -144
right lower quadrant pain | -144
10–15 bowel movements per day | -144
high-grade fever | 0
chills | 0
sweating | 0
tachycardic | 0
heart rate 130 b.p.m. | 0
normotensive | 0
oxygen saturation 94% | 0
posterior oropharynx erythematous | 0
exudates | 0
enlarged cervical lymphadenopathy | 0
tender cervical lymphadenopathy | 0
bilateral cervical lymphadenopathy | 0
left inguinal lymphadenopathy | 0
diffuse abdominal tenderness | 0
scleral injection | 0
mild conjunctivitis | 0
negative SARS-CoV-2 PCR | 0
negative rapid antigen test | 0
leukocytosis | 0
lymphopenia | 0
thrombocytopenia | 0
elevated CRP 27.4 mg/dL | 0
low fibrinogen level 133 mg/dL | 0
D-Dimer 2270 ng/mL FEU | 0
negative blood culture | 0
negative urine culture | 0
negative stool enteric panel | 0
negative respiratory viral panel | 0
right-sided colitis | 0
right mesenteric lymphadenopathy | 0
mild hepatosplenomegaly | 0
normal CXR | 0
started piperacillin–tazobactam | 0
tachycardic | 24
intermittent fevers >102 F | 24
hypotension | 24
IV fluid boluses | 24
transferred to MICU | 24
septic shock | 24
started IV norepinephrine | 24
mild respiratory distress | 24
oxygen saturation 85% | 24
nasal cannula | 24
bilateral pulmonary oedema | 24
elevated pro-BNP >30,000 pg/mL | 24
elevated Troponin T 148.9 ng/L | 24
dilated cardiac chambers | 24
reduced LV systolic function 40–44% | 24
mild global hypokinesis | 24
normal right ventricular systolic function | 24
normal aortic root | 24
small pericardial effusion | 24
mild pulmonic regurgitation | 24
mild tricuspid regurgitation | 24
myocarditis | 24
diagnosed with COVID-19 | -1344
acute colitis | 0
myocarditis | 0
lymphadenopathy | 0
conjunctival injection | 0
negative infectious workup | 0
MIS-C/MIS-A diagnosis | 24
treated with IVIG 2 g/kg | 24
treated with IV methylprednisolone 125 mg | 24
heart rate normalized | 28
defervesced | 28
improvement in abdominal pain | 28
weaned off norepinephrine | 48
transferred out of MICU | 48
IV methylprednisolone transitioned to oral prednisone | 120
heart failure with reduced ejection fraction | 0
started IV furosemide | 0
started angiotensin-converting enzyme inhibitor | 0
discharged on lisinopril | 0
discharged on carvedilol | 0
discharged on furosemide | 0
complete resolution of symptoms | 2160
scheduled for TTE | 2160
