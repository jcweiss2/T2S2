62 years old | 0
female | 0
necrotizing fasciitis of her left thigh and groin | 0
carbuncle | -336
chills | -336
type 2 diabetes mellitus | -6720
ascorbic acid | -6720
hypotensive | 0
blood pressure of 87/63 mm Hg | 0
pulse of 92 bpm | 0
temperature of 36.6°C | 0
severe tenderness to her entire left thigh | 0
posterior crepitus | 0
intravenous fluid resuscitation | 0
hemoglobin of 7.8 g/dl | 0
mean corpuscular volume of 71.9 fl | 0
white blood cell count of 11.9 × 103 µl | 0
platelet count of 151 × 103 µl | 0
reticulocyte count of 3.39% | 0
immature reticulocyte fraction of 35.80% | 0
serum iron level of 7.0 µg/dl | 0
serum transferrin level of 123 mg/dl | 0
total iron-binding capacity of 7.0 µg/dl | 0
direct Coombs test negative | 0
fecal occult blood testing negative | 0
air in the posterior thigh muscles | 0
necrotizing fasciitis | 0
vancomycin | 0
clindamycin | 0
piperacillin/tazobactam | 0
septic shock | 0
fasciotomy | 0
debridement | 0
disarticulation of the left lower extremity | 0
C. septicum | 0
frank blood in her fecal management tube | 288
colonoscopy | 288
fungating polypoid, sessile and ulcerated partially obstructing large mass in her cecum | 288
well-differentiated invasive adenocarcinoma | 288
laparoscopic right hemicolectomy | 297
CT imaging of the abdomen, pelvis, and thorax negative for metastatic spread | 297
no signs or symptoms of recurrence of colon cancer | 8760