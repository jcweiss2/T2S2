25 years old | 0
    woman | 0
    diabetes | 0
    presented to the emergency department | 0
    headache | -168
    right-side neck pain | -168
    shoulder pain | -168
    intermittent fever | -48
    dry cough | -48
    odynophagia | -48
    ill looking | 0
    afebrile | 0
    pulse 115 bpm | 0
    blood pressure 95/60 mm Hg | 0
    respiratory examination normal | 0
    cardiovascular examination normal | 0
    neurological examination normal | 0
    abdominal examination normal | 0
    Kernig's sign negative | 0
    Brudzinski's sign negative | 0
    right-side neck tenderness | 0
    exudative tonsillitis | 0
    WBC count 7.7 | 0
    hemoglobin 10.9 | 0
    thrombocytopenia | 0
    platelet count 22 | 0
    elevated C reactive protein 33.9 | 0
    toxic granulation on blood film | 0
    Na 136 | 0
    K 4.6 | 0
    BUN 14 | 0
    creatinine 0.4 | 0
    AST 27 | 0
    ALT 3 | 0
    direct hyperbilirubinemia | 0
    direct bilirubin 2.0 | 0
    total bilirubin 2.4 | 0
    ECG sinus tachycardia | 0
    initial chest X-ray bilateral infiltrates | 0
    repeat chest X-ray right pleural effusion | 48
    CT neck and chest acute thrombosis right internal jugular vein | 0
    CT septic emboli throughout lung parenchyma | 0
    duplex right upper limb and neck thrombosis right internal jugular vein | 0
    prothrombin 12.7 s | 0
    partial thromboplastin 35.6 s | 0
    INR 1.18 | 0
    HIV negative | 0
    Monospot negative | 0
    Mantoux negative | 0
    antinuclear antibody 1+ fine speckled pattern | 0
    anti-DNA negative | 0
    extractable nuclear antigen panel MI2A++ | 0
    RP11+ | 0
    RP155+ | 0
    C3 157 mg/dL | 0
    C4 26 mg/dL | 0
    cytoplasmic antineutrophil cytoplasmic antibodies negative | 0
    echocardiogram normal | 0
    urine culture no bacterial growth | 120
    blood culture no bacterial growth | 120
    commenced ceftriaxone | 0
    day 2 post hospitalization | 48
    markedly distressed | 48
    acidotic pH 7.159 | 48
    transferred to ICU | 48
    ventilatory support | 48
    meropenem | 48
    vancomycin | 48
    vasopressors | 48
    anticoagulated with rivaroxaban | 48
    acute kidney injury | 48
    creatinine rise to 1.9 mg/dL | 48
    creatinine resolved | 432
    full recovery | 480
    discharged | 480
    oral anticoagulants | 480
    oral antibiotics | 480
    insulin therapy | 480
    scheduled follow-up outpatient medical clinic | 480
    scheduled follow-up diabetes clinic | 480
    acute tonsillitis | 0
    thrombophlebitis | 0
    internal jugular vein thrombosis | 0
    septic emboli to lungs | 0
    Lemierre's syndrome | 0
    neck pain | 0
    fever | 0
    dry cough | 0
    odynophagia | 0
    sore throat | -168
    swollen neck | 0
    tender neck | 0
    deranged liver enzymes | 0
    hyperbilirubinemia | 0
    acute viral pharyngitis | 0
    negative blood cultures | 120
    F. necrophorum | 0
    necrotic abscesses | 0
    thrombosis internal jugular vein | 0
    septic emboli lungs | 0
    oropharyngeal sepsis | 0
    metastatic infection | 0
    viral pharyngitis | 0
    pneumonia | 0
    infective endocarditis | 0
    acute retroviral illness | 0
    infectious mononucleosis | 0
    leptospirosis | 0
    ceftriaxone | 0
    meropenem | 48
    vancomycin | 48
    acute respiratory distress | 48
    ventilation | 48
    clindamycin | 0
    cefoxitin | 0
    imipenem | 0
    metronidazole | 0
    penicillin | 0
    macrolides resistant | 0
    gentamicin resistant | 0
    quinolones resistant | 0
    acute respiratory distress syndrome | 48
    improvement after 5 days ICU | 120
    managed in medical ward | 120
    anticoagulation therapy | 48
    surgical management ligation/resection internal jugular vein | 0
    persistent septic embolization | 0
    acute renal failure | 48
    resolved with fluids and antibiotics | 432
    bone and joint complications | 0
    septic arthritis | 0
    osteomyelitis | 0
    skin and soft tissue lesions | 0
    purulent meningitis | 0
    endocarditis | 0
    pericarditis | 0
    <|eot_id|>
    