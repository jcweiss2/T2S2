55 years old | 0  
    female | 0  
    non-insulin dependent diabetes | 0  
    midline lower abdominal pain | -96  
    dysuria | -96  
    lower back pain | -96  
    nausea | -96  
    vomiting | -96  
    vaginal bleeding | -96  
    amenorrhea | -2880  
    afebrile | 0  
    normotensive | 0  
    non-tachycardic | 0  
    normal cardiovascular exam | 0  
    general lower abdominal tenderness | 0  
    enlarged uterus | 0  
    pelvic exam | 0  
    normal external female genitalia | 0  
    displaced cervix anteriorly | 0  
    no cervical motion tenderness | 0  
    cervix not directly visualized | 0  
    wet prep negative | 0  
    endometrial biopsy | 0  
    leukocytosis (19 k/mm3) | 0  
    urinalysis with nitrites | 0  
    urinalysis with leukocytes | 0  
    urinalysis with blood | 0  
    urinalysis with leukocytosis | 0  
    transvaginal ultrasound showing uterine masses | 0  
    leiomyomata | 0  
    largest fibroid fundal (6 cm) | 0  
    fibroids affecting endometrium and serosa | 0  
    thickened endometrium (46.9 mm) | 0  
    lobulated tissue in cavity | 0  
    ovaries not visualized | 0  
    acute cystitis | 0  
    degenerating fibroids | 0  
    underlying malignancy | 0  
    pain improved with acetaminophen | 0  
    pain improved with ibuprofen | 0  
    treated for acute cystitis | 0  
    discharged home | 0  
    worsening suprapubic pain | 96  
    fevers | 96  
    chills | 96  
    nausea | 96  
    vomiting | 96  
    vaginal bleeding | 96  
    no malodorous discharge | 96  
    lower abdominal tenderness | 96  
    suprapubic tenderness | 96  
    pelvic exam unchanged | 96  
    initially afebrile | 96  
    normal heart rate | 96  
    hypotensive (systolic 60-90) | 96  
    hypotensive (diastolic 30-50) | 96  
    leukocytosis (17 k/mm3) | 96  
    elevated lactate (4.0 mmol/L) | 96  
    CT abdomen and pelvis findings | 96  
    fibroid uterus | 96  
    pelvic free fluid | 96  
    expanded endometrial cavity (8 cm) | 96  
    hyperdensity (4 cm) | 96  
    sepsis due to urinary source | 96  
    gynecologic source | 96  
    gastrointestinal source | 96  
    crystalloid fluid resuscitation | 96  
    norepinephrine started | 96  
    broad spectrum antibiotics (vancomycin, piperacillin-tazobactam) | 96  
    admitted to MICU | 96  
    leukocytosis improved (9.5 k/mm3) | 96  
    lactate improved (3.6 mmol/L) | 96  
    persistent hypotension | 96  
    mild tachycardia | 96  
    afebrile | 96  
    serial physical exams | 96  
    serial laboratory exams | 96  
    antibiotics continued | 96  
    worsening leukocytosis (66.3 k/mm3) | 105  
    lactic acidosis (4.9 mmol) | 105  
    required vasopressin | 105  
    antibiotics broadened to meropenem | 105  
    minimal urine output (220 ml) | 105  
    lower abdominal guarding | 105  
    exploratory laparotomy | 105  
    total abdominal hysterectomy | 105  
    bilateral salpingo-oophorectomy | 105  
    pressor support required | 105  
    enlarged uterus (20 cm) | 105  
    necrotic intrauterine mass (8 cm) | 105  
    foul-smelling mass | 105  
    no myometrial invasion | 105  
    uncomplicated surgery | 105  
    estimated blood loss (150 ml) | 105  
    abdomen irrigated with saline | 105  
    Blake drain placed | 105  
    fascia closed | 105  
    subcutaneous tissue packed | 105  
    pressor support decreased | 105  
    urine output increased | 105  
    extubated | 105  
    transferred to SICU | 105  
    weaned off vasopressors | 120  
    blood cultures: Clostridium species | 120  
    blood cultures: Bacteroides vulgatus | 120  
    antibiotics narrowed (ampicillin-sulbactam, clindamycin) | 120  
    transferred out of SICU | 168  
    post-operative milestones met | 168  
    IV antibiotics continued | 288  
    white blood cell count normalized | 288  
    discharged home | 288  
    wound-vac | 288  
    amoxicillin-clavulanate | 288  
    metronidazole | 288  
    surgical pathology: pT1a carcinosarcoma | 288  
    adjuvant carboplatin | 288  
    adjuvant paclitaxel | 288  
    vaginal brachytherapy | 288  
    
