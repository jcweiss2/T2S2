30 years old | 0
female | 0
abdominal pain | -48
nausea | -48
vomiting | -48
fever | -48
severe pulmonary hypertension | 0
bilateral pulmonary emboli | 0
right heart failure | 0
hypothyroidism | 0
systemic hypertension | 0
WHO functional class III | 0
tenderness to palpation over the right lower quadrant | 0
leukocytosis | 0
left shift | 0
CT scan of the abdomen and pelvis | 0
distended fluid-filled appendix | 0
appendicoliths | 0
surrounding edema | 0
respiratory distress | 0
admitted to the intensive care unit | 0
right heart catheterization | 0
severe pulmonary hypertension | 0
right ventricular systolic pressure of 120 mm Hg | 0
moderate to severe tricuspid regurgitation | 0
sildenafil | 0
intravenous epoprostenol | 0
heparin infusion | 0
intravenous piperacillin/tazobactam | 0
worsening leukocytosis | 24
fever of 39.1°C | 24
tachypnea | 24
worsening focal peritonitis | 24
severe sepsis | 24
impending shock | 24
femoral vessel cannulation | 24
open appendectomy | 24
purulent peritoneal fluid | 24
necrotic and gangrenous appendix | 24
multiple perforations | 24
abdominal cavity irrigation | 24
abdomen closed with a Jackson-Pratt drain | 24
extubated | 24
transferred to the intensive care unit | 24
arterial and venous sheaths removed | 48
discharged | 432
postoperative day 18 | 432
sildenafil | 432
bumetanide | 432
macitentan | 432
intravenous epoprostenol | 432