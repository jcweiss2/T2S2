27 years old | 0
male | 0
admitted to the hospital | 0
abdominal pain | -24
vomiting | -24
blunt abdominal trauma | -24
high heart rate | 0
respiratory rate | 0
blood pressure | 0
temperature | 0
oxygen saturation level | 0
generalized abdominal pain | 0
voluntary muscular defense | 0
signs of peritoneal irritation | 0
normal hemoglobin level | 0
mild leukocytosis | 0
rupture of the third portion of the duodenum | 0
retropneumoperitoneum | 0
exploratory laparotomy | 0.5
free perforation | 0.5
duodenorrhaphy | 1
Connel-Mayo suture | 1
Lambert suture | 1
vascular prolene | 1
Jackson-Pratt drain | 1
nasogastric tube | 1
piperacillin-tazobactam antibiotic | 1
enteral nutrition | 1
peritoneal fluid culture | 24
Enterobacter cloacae complex | 24
inducible strain | 24
beta-lactamases | 24
AmpC pattern | 24
ertapenem | 48
discharged | 168
postoperative control | 168
early diet | 168
physical therapy | 168
early mobilization | 168
restricted sports activity | 168
hospitalization | 0
antibiotic treatment | 1
secondary peritonitis | 1
uncontained perforation | 0
infectology service | 24
elevated acute phase reactants | 24
leukocytosis | 24 
drain removed | 360 
no complications | 720 
no affectation in activities of daily living | 720