female | 0
infant | 0
born via spontaneous vaginal delivery | 0
gestational age of 36 weeks and 0 days | 0
birth weight was 2356 g | 0
Apgar scores were 9 at both 1 and 5 minutes | 0
meconium staining was not observed | 0
preterm premature rupture of membranes | -168
prescribed intravenous ampicillin | -168
cultures of vaginal and stool samples were positive for Group B Streptococcus | -336
respiratory distress | 0
resuscitation with positive pressure ventilation | 0
admitted to the neonatal intensive care unit | 0
placed on a mechanical ventilator | 0
work-up for sepsis | 0
blood cultures | 0
antibiotics were not administered | 0
fever | 16
convulsions | 16
drowsiness | 16
pale | 16
cold extremities | 16
cyanosis of the extremities | 16
poor capillary refill | 16
body temperature of 38.8 °C | 16
pulse of 170 beats per minute | 16
blood pressure of 60/35 mmHg | 16
respiratory rate of 80 breaths per minute | 16
oxygen saturation of 87% on mechanical ventilation | 16
cardiovascular examination was normal | 16
lungs were clear on auscultation | 16
abdomen was soft | 16
muscle tone was slightly increased | 16
no evidence of a skin rash | 16
no subcutaneous hemorrhage | 16
diagnostic assessment | 16
laboratory findings consistent with disseminated intravascular coagulation | 16
cerebrospinal fluid examination | 16
high cell count | 16
glucose concentration of 0.06 mmol/L | 16
gram-negative rod organisms | 16
abdominal US performed | 16
bilateral adrenal hemorrhage | 16
Waterhouse-Friderichsen syndrome | 16
central diabetes insipidus | 72
lethargy | 72
blood pressure decreased to 50/30 mmHg | 72
urine output increased to 10 mL/kg per hour | 72
urine had a specific gravity of 1.005 | 72
osmolality of 160 mOsm/kg H2O | 72
serum sodium concentration of 155 mmol/L | 72
serum osmolality of 332 mOsm/kg H2O | 72
serum antidiuretic hormone level of 1.3 pg/mL | 72
treated with appropriate antibiotics | 16
hydrocortisone | 16
blood pressure returned to the normal range | 40
no further steroid therapy | 72
follow-up examinations showing a gradual regression of AH | 72
blood and CSF cultures after 36 hours of treatment were both negative | 52
treatment with antibiotics was continued | 16
treated with intravenous vasopressin | 96
urine output decreased to 4 mL/kg/h | 120
urine osmolality improved to 213 mOsm/kg H2O | 120
vasopressin dose was reduced | 120
intravenous vasopressin was discontinued | 288
cerebral magnetic resonance imaging | 240
bilateral encephalomalacia | 240
minor bleeding | 240
splenial lesion | 240
mild encephalitis/encephalopathy | 240
reversible splenial lesion | 240
no signs of abscess | 240
no ventriculitis | 240
no pituitary gland abnormality | 240
endocrine assessments | 840
serum concentrations of thyroid-stimulating hormone | 840
thyroid hormone | 840
adrenocorticotropic hormone | 840
early morning cortisol level was low | 840
corticotropin-releasing hormone stimulation test | 840
normal adrenocorticotropic hormone response | 840
no evidence of central adrenal insufficiency | 840
automated auditory brainstem response testing | 840
electroencephalography | 840
no abnormalities | 840
discharged | 1080