37 years old| 0
    pregnant woman (G3P2)| 0
    presented to the emergency department| 0
    33 weeks' gestation| 0
    breathlessness| -216
    tested positive for COVID-19| -216
    feeling generally unwell| -216
    non-productive cough| -216
    took to her bed| -216
    little oral intake| -216
    little fluid intake| -216
    increase in work of breathing| -72
    unable to mobilise short distances| -72
    denied chest pain| 0
    denied calf tenderness| 0
    denied orthopnoea| 0
    denied paroxysmal nocturnal dyspnoea| 0
    well-controlled asthma| 0
    gastric sleeve surgery| 0
    regular inhalers| 0
    vitamin B12 injections| 0
    non-smoker| 0
    no regular alcohol| 0
    no illicit medications| 0
    no over-the-counter medications| 0
    hyperemesis gravidarum in the first trimester| -1848
    respiratory rate 32 breaths/min| 0
    oxygen saturations 95% on 4 L/min inspired oxygen| 0
    heart rate 105 beats/minute| 0
    blood pressure 100/60 mmHg| 0
    apyrexial| 0
    breathless at rest| 0
    Kussmaul breathing| 0
    ketotic breath| 0
    unable to complete full sentences| 0
    bi-basal crepitations| 0
    no wheeze| 0
    clinically dehydrated| 0
    normal neurological examination| 0
    normal cardiovascular examination| 0
    normal abdominal examination| 0
    normal oral glucose tolerance test| 0
    normal glycated haemoglobin A1c| 0
    sinus tachycardia| 0
    chest X-ray confirmed COVID-19 pneumonitis| 0
    CT pulmonary angiography confirmed COVID-19 pneumonitis| 0
    no pulmonary emboli| 0
    metabolic acidosis| 0
    normal blood glucose levels| 0
    normal lactate levels| 0
    denial of toxin ingestion| 0
    denial of drug abuse| 0
    denial of alcohol abuse| 0
    normal renal function| 0
    elevated ketones| 0
    high anion gap| 0
    severe COVID9 infection| 0
    starvation ketosis of pregnancy| 0
    history of gastric bypass surgery| 0
    history of hyperemesis gravidarum| 0
    chronic starvation| 0
    anorexia while acutely unwell| 0
    MDT discussion| 0
    initiation of treatment for COVID9| 0
    initiation of treatment for metabolic disturbance| 0
    oxygen to maintain saturations >94%| 0
    intramuscular dexamethasone for fetal lung maturity| 0
    prednisolone initiated| 0
    tocilizumab initiated| 0
    administration of corticosteroids discussed| 0
    intravenous 20% dextrose| 0
    intravenous 0.9% sodium chloride| 0
    intravenous 1.6% bicarbonate| 0
    variable rate insulin infusion| 0
    potassium replacement| 0
    Pabrinex| 0
    resolution of metabolic ketoacidosis over 24 hours| 24
    respiratory rate 26 breaths/min| 24
    oxygen saturations 96% on 4 L/min inspired oxygen| 24
    heart rate 100 beats/min| 24
    blood pressure 110/64 mmHg| 24
    apyrexial| 24
    stopped intravenous 20% dextrose| 24
    stopped intravenous 0.9% sodium chloride| 24
    stopped intravenous 1.6% bicarbonate| 24
    stopped variable rate insulin infusion| 24
    stopped potassium replacement| 24
    stopped Pabrinex| 24
    continued prednisolone| 24
    added low molecular weight heparin| 24
    venous thromboembolism prophylaxis| 24
    remained stable over next 6 days| 168
    oxygen saturations deteriorated to 88%| 168
    worsening pneumonitis| 168
    pneumomediastinum| 168
    right apical pneumothorax| 168
    MDT discussion| 168
    decision to deliver the baby| 168
    commenced on ECMO| 168
    delivery| 168
    baby admitted to special care baby unit| 168
    good recovery of baby| 168
    decannulated from ECMO| 408
    discharged from hospital| 408
    well at follow-up 3 months later| 2160
    <|eot_id|>