65 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
admitted to the hospital | 0 | 0 | Factual
fever | 0 | 48 | Factual
chills | 0 | 48 | Factual
pain in left leg | 0 | 48 | Factual
parkinsonism | -8760 | 0 | Factual
diabetes mellitus | -8760 | 0 | Factual
levodopa / carbidopa | -8760 | 0 | Factual
rasagiline | -8760 | 48 | Factual
ropinirole | -8760 | 0 | Factual
trihexyphenidyl | -8760 | 0 | Factual
amantadine | -8760 | 0 | Factual
metformin | -8760 | 48 | Factual
glipizide | -8760 | 48 | Factual
cellulitis | 0 | 48 | Factual
intravenous clindamycin | 0 | 48 | Factual
intravenous benzylpenicillin | 0 | 48 | Factual
high-temperature spikes | 72 | 72 | Factual
tachycardia | 72 | 72 | Factual
tachypnea | 72 | 72 | Factual
hypotensive | 72 | 72 | Factual
encephalopathic | 72 | 72 | Factual
shifted to ICU | 72 | 72 | Factual
intravenous linezolid | 72 | 120 | Factual
intravenous piperacillin with tazobactam | 72 | 120 | Factual
vancomycin not considered | 72 | 72 | Factual
hemodynamics improved | 72 | 120 | Factual
minimal inotropic supports | 72 | 120 | Factual
oral hypoglycemic agents stopped | 72 | 72 | Factual
switched to insulin | 72 | 120 | Factual
confused | 96 | 120 | Factual
drowsy | 96 | 120 | Factual
disoriented | 96 | 120 | Factual
altered sensorium | 96 | 120 | Factual
myoclonus | 96 | 120 | Factual
tremors | 96 | 120 | Factual
jerky movements | 96 | 120 | Factual
no neck stiffness | 96 | 120 | Factual
computed tomography of the brain | 96 | 96 | Factual
cerebrospinal fluid analysis | 96 | 96 | Factual
improving white blood cell counts | 96 | 120 | Factual
better glycemic control | 96 | 120 | Factual
sterile blood and pus cultures | 96 | 120 | Factual
serotonin syndrome suspected | 120 | 120 | Factual
linezolid stopped | 120 | 120 | Factual
rasagiline stopped | 120 | 120 | Factual
temperature settled | 128 | 128 | Factual
heart rate normal | 144 | 144 | Factual
sensorium improved | 144 | 144 | Factual
tremors subsided | 144 | 144 | Factual
shifted out of ICU | 192 | 192 | Factual
started walking with support | 240 | 240 | Factual
discharged from the hospital | 240 | 240 | Factual
anti-parkinsonism drugs | 240 | 0 | Factual
rasagiline added | 240 | 0 | Factual
regular follow-up with neurologist | 240 | 0 | Factual
stable and asymptomatic for serotonin syndrome | 240 | 0 | Factual