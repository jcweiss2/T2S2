48 years old | 0
male | 0
SARS-CoV-2 infection | -168
ground-glass pattern on thoracic computed tomography | -168
positive nasopharyngeal swab test | -168
oseltamivir | -168
hydroxychloroquine | -168
broad-spectrum antibiotics | -168
endotracheal intubation | -144
invasive mechanical ventilation | -144
favipiravir | -144
ARDS | -144
rehabilitation program | -144
in-bed positioning | -144
passive range of motion | -144
prone position | -144
cytokine storm syndrome | -72
candidemia | -72
intravenous tocilizumab | -72
immune plasma | -72
intravenous high-dose glucocorticoids | -72
antifungal therapy | -72
controlled breathing techniques | 0
bronchial hygiene-airway clearance techniques | 0
home-based respiratory muscle exercise program | 0
threshold inspiratory muscle trainer | 0
admitted to the inpatient clinic of the Department of Physical Medicine and Rehabilitation | 0
weakness | 0
distal muscles of the upper and lower extremities | 0
right wrist drop | 0
bilateral foot drop | 0
symmetrical mild distal muscle atrophy | 0
contractures of the left hip and left knee | 0
sacral decubitus ulcer | 0
sensorimotor axonal peripheral neuropathy | 0
ICU-AW | 0
rehabilitation program | 0
Mini-Mental State Examination | 0
General Health Perception | 0
Mental Health Perception | 0
Physical Function | 0
functional ambulation category | 0
muscle strength score | 0
postural hypotensive attacks | 0
tilt table | 0
active-assisted and active ROM | 0
isometric strength exercises | 0
isotonic strength exercises | 0
mobilization | 0
methenolone enanthate | 0
neuromuscular electrical stimulation | 0
collagen-containing dressing | 0
high-density ankle-foot orthosis | 0
walker | 0
improved cognitive scores | 168
improved quality of life | 168
improved life activity scales | 168
discharge | 168
MMSE | 168
General Health Perception | 168
Mental Health Perception | 168
Physical Function | 168
muscle strength | 168
fine motor grip skills | 168
hand grip strength | 168
pinch strength | 168