56 years old | 0
woman | 0
presented to a community hospital | 0
weakness | -720
numbness | -720
weakness in lower extremities | -720
numbness and weakness in lower extremities | -720
numbness and weakness in lower extremities progressing to hands and neck | -720
numbness and weakness in lower extremities progressing to hands and neck over a few days | -720
type 2 diabetes mellitus | -17520
hypertension | -17520
episode of necrotizing pancreatitis due to gallstones | -17520
severe protein-calorie malnutrition | -17520
total parenteral nutrition | -17520
discontinued total parenteral nutrition | -4320
returned to a normal diet | -4320
lumbar puncture | 0
albuminocytologic dissociation in cerebrospinal fluid | 0
presumptive diagnosis of Guillain-Barré syndrome | 0
presumptive diagnosis of acute inflammatory demyelinating polyradiculoneuropathy | 0
brain MRI scan showing small vessel ischemic changes | 0
empiric intravenous immunoglobulin treatment | 0
no clinical response | 120
worsening pancytopenia | 120
encephalopathy | 120
transfer to a specialist center | 120
hypotensive | 0
blood pressure 64/48 mmHg | 0
unresponsive to verbal stimuli | 0
minimally responsive to painful stimuli | 0
Glasgow Coma Scale score of 6 | 0
anasarcic | 0
flaccid paralysis of all four extremities | 0
calcium 6.7 mg/dL | 0
hemoglobin 9.4 g/dL | 0
white cell count 2.1×10^9/L | 0
phosphorus 1.1 mg/dL | 0
creatinine <0.2 mg/dL |#generated by assistant
albumin <1.5 gm/dL | 0
lactate 4 mmol/L | 0
nutritional risk screening score 5 | 0
malnutrition universal screening score 5 | 0
intubation | 0
resuscitated with intravenous fluids | 0
required intravenous infusion of norepinephrine | 0
meropenem treatment | 0
vancomycin treatment | 0
anidulafungin treatment | 0
provisional diagnosis of AIDP complicated by septic shock | 0
empirical treatment with high-dose intravenous thiamine | 0
electroencephalogram showing diffuse slow waves | 0
no seizure activity | 72
brain MRI scan showing hyperintensity of bilateral medial thalamus | 72
serum thiamine level 104 nmol/L | 72
mental status markedly improved | 96
able to understand simple commands | 96
norepinephrine discontinued | 96
antimicrobial treatment discontinued | 96
resolution of hemodynamic stability | 96
negative blood cultures | 96
negative urine cultures | 96
successfully extubated | 120
electromyography showing severe sensorimotor polyneuropathy | 168
mentation improved | 168
weakness improved | 168
transferred out of ICU | 336
thiamine supplementation continued | 336
discharged | 336
