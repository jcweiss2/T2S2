32 years old | 0
    male | 0
    presented to emergency department | 0
    painful right lower limb swelling | -120
    difficulty to walk | -120
    generalized weakness | -120
    fever | -120
    hepatitis C | 0
    intravenous drug abuse | 0
    last use 5 days ago | -120
    groin region | -120
    focal tenderness | 0
    ecchymosis | 0
    marked edema of knee joint | 0
    admitted to department of pathology | 0
    synovial fluid aspiration | 0
    synovial fluid culture sent | 0
    neurological examination satisfactory | 0
    vascular examination satisfactory | 0
    cellulitis diagnosis | 0
    septic arthritis suspicion | 0
    piperacillin administration | 0
    metronidazole administration | 0
    intravenous fluids | 0
    blood pressure 98/54 mmHg | 0
    heart rate 123 b/min | 0
    respiratory rate 22/min | 0
    oxygen saturation 92% | 0
    temperature 38.1°C | 0
    alert | 0
    oriented | 0
    neurovascularly intact | 0
    nonsteroidal anti-inflammatory drugs | 0
    white blood cells 11,060/μL | 0
    C-reactive protein 36.8 mg/dL |9
    hematocrit 40.7% | 0
    hemoglobin 14.3 g/dL | 0
    platelets 184,000/μL | 0
    D-dimers 127,5 μg/L | 0
    urea 100 mg/dL | 0
    creatinine 0.81 mg/dL | 0
    erythrocyte sedimentation rate 108 mm/h | 0
    Na 145 mmol/L | 0
    K 4.6 mmol/L | 0
    creatine kinase 1210 IU/L | 0
    lactate dehydrogenase 355 IU/L | 0
    cutaneous ecchymosis worsened | 0
    contrast-enhanced CT scan | 0
    inflammatory stranding | 0
    low attenuation | 0
    necrosis suspicion in rectus femoris | 0
    necrosis suspicion in vastus lateralis | 0
    NF suspicion | 0
    knee arthrotomy | 0
    extensive synovectomy | 0
    irrigation with 9 L saline | 0
    debridement of infected soft tissues | 0
    fasciotomy through anterolateral approach | 0
    debridement of subcutaneous fat necrosis | 0
    debridement of vastus lateralis necrosis | 0
    S. aureus infection confirmation | 0
    vancomycin addition | 0
    ICU admission | 0
    daily wound evaluation | 24
    irrigation | 24
    aggressive surgical debridement | 24
    lesions worsened | 168
    foul-smelling necrotic materials | 168
    surgical exploration | 168
    necrosis removal | 168
    major vessel bleeding | 168
    angiography | 168
    popliteal artery thrombosed aneurysm | 168
    peroneal artery thrombosed aneurysm | 168
    hematoma/thrombus evacuation | 168
    stent insertion | 168
    clinical condition improved | 480
    reconstructive surgery scheduled | 480
    plastic surgery scheduled | 480
    clinical picture deteriorated | 720
    septic shock | 720
    above-the-knee amputation | 720
    ICU stay | 720
    metabolic support | 720
    hemodynamic support | 720
    transferred to department | 2496
    local wound care | 2496
    fluid management | 2496
    discharge | 4176
    follow-up | 4176
    