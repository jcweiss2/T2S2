48 years old | 0
male | 0
admitted to urology | 0
necrotic lesion on glans penis | 0
sepsis | 0
infected calciphylaxis-related ulcer on thigh | 0
broad spectrum antibiotics | 0
increasing bladder volumes | 0
urinary tract infection | 0
infrequent episodes of urinary incontinence | -672
end-stage renal failure | -672
peritoneal dialysis | -672
haemodialysis | -1344
calciphylaxis | -1344
type 2 diabetes | -672
cerebrovascular accident | -672
atrial fibrillation | -672
palpable bladder | 0
tender necrotic lesion | 0
ultrasound scan | -336
bladder scan | 0
ultrasound guided aspiration of bladder | 0
apixaban | 0
protracted admission | 24
slow resolution of infected ulcer | 24
physical deconditioning | 24
further aspiration of bladder | 2160
stable lesion | 2160
discharged to nursing home | 4320
urinary diversion | 4320
suprapubic catheter | 4320
urinary retention | 0
meatal obstruction | 0
painless retention | 0
catheter-associated UTI | 0
sepsis due to UTI | 0
aspiration on triannual basis | 4320
calciphylaxis diagnosis | -1344
poor prognosis | -1344
yearly mortality | -1344
punch biopsy | -1344
wound care | 0
analgesia | 0
infection prevention | 0
treatment | 0
regulation of serum vitamin D | 0
regulation of serum calcium | 0
regulation of serum phosphate | 0
diet modification | 0
calcium and phosphate chelating agents | 0
Cinacalcet | 0
sodium thiosulfate | 0
haemodialysis | 0
surgical intervention | 0
debridement | 0
partial penectomy | 0
total penectomy | 0
urinary diversion | 0
parathyroidectomy | 0
hyperparathyroidism | -1344
penile calciphylaxis | -1344
necrotic lesions | -1344
vascular calcification | -1344
thrombosis formation | -1344
radiological investigations | 0
ultrasound | 0
CT | 0
MRI | 0
urinary retention with meatal obstruction | -672
suprapubic catheter insertion | -672
patient satisfaction | -672
surgical debridement | -672
temporary urethral catheters | -672
total penectomy | -672
perineal urethrostomy formation | -672
nosocomial UTI | 0
catheterisation | 0
UTI risk | 0
sepsis risk | 0
mortality risk | 0
aspiration on triannual basis | 4320
low risk management option | 4320
obstructed urinary tract | 0
life expectancy | -1344
reduced physiological reserves | -1344
sepsis secondary to catheter associated UTI | 0
fatal outcome | 0
interval sterile ultrasound guided aspiration | 4320
safer method of bladder management | 4320