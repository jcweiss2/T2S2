73 years old | 0
female | 0
fever | -168
asthenia | -168
odynophagia | -168
epistaxis | -168
cacosmia | -2628
foul-smelling nasal crusts | -2628
diabetes | 0
hypertension | 0
admitted to the hospital | 0
afebrile | 0
oriented | 0
cooperative | 0
crackles in the lung bases | 0
mucopurulent secretion in the left external auditory canal | 0
peritonsillar bulging | 0
hyperemia | 0
intravenous antibiotic therapy with ceftriaxone and clindamycin | 0
puncture of the oral bulge | 24
no secretion was drained | 24
second puncture | 48
larvae coming out through the mouth and left nostril | 48
septicemia | 72
decreased level of consciousness | 72
blood desaturation | 72
intubation | 72
mechanical ventilation | 72
iodoform applied to the oral cavity and nasal passages | 72
ivermectin administered | 72
piperacillin/tazobactam and vancomycin administered | 72
otorhinolaryngological examination | 72
removal of larvae | 72
computed tomography of the nose and paranasal sinuses | 96
computed tomography of the temporal bones, skull, and lung | 96
complete removal of larvae | 120
respiratory failure | 720
pneumonia | 720
death | 720