77 years old | 0
male | 0
admitted to the hospital | 0
abrupt onset of impaired consciousness | 0
hypotension | 0
intermittent mild lower abdominal discomfort | -120
bloody loose stools | -120
prostate cancer | -8760
Bicalutamide | -8760
hypertension | 0
hyperlipidemia | 0
hyperuricemia | 0
lumbar spinal stenosis | 0
Glasgow score 10 | 0
limbs were cold and moist | 0
body temperature 35.6 °C | 0
pulse rate 42 bpm | 0
blood pressure 65/36 mmHg | 0
respiration rate 28 breaths/min | 0
oxygen saturation 95 % | 0
mild abdominal distension | 0
normal bowel sounds | 0
normal white blood cell count | 0
normal platelet count | 0
normal hemoglobin level | 0
elevated serum creatinine | 0
elevated lactic acid | 0
elevated hemoglobin A1c | 0
echocardiography demonstrated no abnormalities | 0
abdominal ultrasound demonstrated no abnormalities | 0
non-contrast-enhanced whole-body CT revealed mild edematous swelling of the small-intestinal wall | 0
septic shock | 0
intravenous crystalloid solution administered | 0
noradrenaline administered | 0
Meropenem initiated | 0
state of consciousness improved | 72
vital signs normalized | 72
spike in body temperature | 72
C. paraputrificum grown from blood culture | 0
ampicillin/sulbactam treatment | 0
laboratory parameters improved | 96
clinical conditions improved | 96
discharged from ICU | 96
abdominal manifestations persisted | 96
low-grade fever | 96
mild anemia | 96
Clostridium difficile toxins A and B negative | 96
glutamate dehydrogenase antigen negative | 96
stools negative for ova, parasites, and culture | 96
sigmoidoscopy demonstrated diffuse mucosal inflammation | 840
histopathology revealed crypt disarray | 840
ulcerative colitis diagnosed | 840
oral probiotics administered | 840
intestinal prokinetic medications administered | 840
abdominal X-ray demonstrated dilated colon | 1488
non-contrast-enhanced abdominal CT confirmed colonic dilatation | 1488
ACPO diagnosed | 1488
total parenteral nutrition initiated | 1488
pharmacologic and endoscopic decompression therapy initiated | 1488
dilated colon resected | 2232
C. paraputrificum bacteremia | 0
und diagnosed ulcerative colitis | 0
acute colonic pseudo-obstruction | 1488