left lower quadrant abdominal pain | -168
pelvic heaviness | -168
urinary frequency | -168
miscarriages | -10080
tubal ligation | -10080
active smoker | 0
no medication | 0
large and painful mass | 0
pelvic MRI | 0
mass measuring 18 × 17 × 12 cm | 0
no lymphadenopathy | 0
no ascites | 0
no peritoneal implants | 0
normal uterus and adnexa | 0
negative serum tumor markers | 0
surgical pelvic exploration | -744
mass of the left broad ligament | -744
no ascites | -744
no peritoneal carcinomatosis | -744
normal uterus and right adnexa | -744
total hysterectomy with adnexectomy | -744
removal of the mass | -744
definitive histological diagnosis of leiomyosarcoma | -744
isolated fever | 48
major inflammatory syndrome | 48
leukocytes 15,000/μL | 48
C-reactive protein 317 mg/dL | 48
contrast-enhanced computed tomography scan | 48
abscess | 48
blood pressure dropped | 48
intravenous volume replacement with 2 L of Ringer Lactate | 48
vasopressor therapy | 48
emergency revision surgery | 48
peritoneal cavity exploration | 48
moderately abundant non-purulent serosanginous peritoneal fluid | 48
adhesions to the Douglas pouch | 48
peritonitis | 48
antibacterial treatment with piperacillin/tazobactam and gentamicin | 48
extubation | 72
hemodynamic support with noradrenaline | 72
decrease in noradrenaline requirement | 96
discontinuation of noradrenaline | 96
decrease in inflammatory markers | 96
microbiological analysis of the peritoneal fluid | 96
identification of Gardnerella vaginalis | 96
discontinuation of gentamicin | 96
addition of metronidazole | 96
identification of Atopobium vaginae | 120
sterile preoperative blood cultures | 120
antibacterial susceptibility testing of Gardnerella vaginalis | 120
antibacterial susceptibility testing of Atopobium vaginae | 120
discharge from intensive care unit | 120
stop of antibacterial therapy | 168