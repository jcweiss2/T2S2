14 years old | 0 | 0 
male | 0 | 0 
admitted to the hospital | 0 | 0 
near-drowning incident | -1 | -1 
cardiopulmonary resuscitation (CPR) | -1 | -1 
abdominal pain | 0 | 0 
diffuse abrasions on torso | 0 | 0 
pneumoperitoneum | 0 | 0 
pneumomediastinum | 0 | 0 
intraabdominal free fluid | 0 | 0 
taken to the operating room | 0 | 0 
gross contamination with food debris | 0 | 0 
total gastroesophageal junction (GEJ) disruption | 0 | 0 
patient became hemodynamically labile | 0 | 0 
damage control procedure | 0 | 0 
distal esophagus and proximal stomach stapled closed | 0 | 0 
four drains placed | 0 | 0 
gastrostomy (G) tube placed | 0 | 0 
mediastinal drain placed | 0 | 0 
large bore nasogastric (NG) tube placed | 0 | 0 
fascia closed | 0 | 0 
transferred to Pediatric Intensive Care Unit (ICU) | 0 | 0 
septic shock | 0 | 18 
respiratory failure | 0 | 18 
prolonged intubation | 0 | 18 
deep venous thrombosis | 0 | 18 
pulmonary embolism | 0 | 18 
bilateral pleural effusions | 0 | 18 
general deconditioning | 0 | 18 
parenteral nutrition started | 0 | 18 
extubated | 18 | 18 
fluoroscopic evaluation | 18 | 18 
leak in esophagus | 18 | 18 
stomach negative for leak | 18 | 18 
enteral nutrition initiated via G tube | 18 | 18 
discharged | 50 | 50 
nasogastric tube and mediastinal drain | 50 | 120 
Ivor-Lewis distal esophagectomy | 120 | 120 
gastric pull-up for esophagogastric anastomosis | 120 | 120 
gastric conduit made | 120 | 120 
right thoracotomy performed | 120 | 120 
distal esophagus identified | 120 | 120 
tubularized portion of stomach advanced into chest | 120 | 120 
esophagogastric anastomosis | 120 | 120 
leak test performed | 120 | 120 
jejunostomy tube placed | 120 | 120 
extubated | 123 | 123 
nutritionally supported with jejunostomy enteral feeds | 123 | 130 
esophagram showed no leak | 130 | 130 
initiated on liquid diet | 130 | 130 
discharged | 130 | 130 
tolerate regular diet | 155 | 155 
gaining weight and recovering well | 155 | 155