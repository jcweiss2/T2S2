64 years old | 0
female | 0
diabetes mellitus | -8760
admitted to the intensive care unit | 0
septic shock | 0
acute left pyelonephritis | 0
CT scan | 0
lower mass syndrome of the left kidney | 0
necrosis | 0
calcifications | 0
wide nephrectomy with adrenalectomy | 24
kidney occupied at its inferior pole by a fleshy well-defined tumor | 24
tumor measuring 7.5 × 7 × 7 cm | 24
solid on cutting with patchy hemorrhagic and necrotic areas | 24
dual carcinomatous proliferation composed of clear and eosinophilic cells | 24
lobular growth pattern | 24
tubulo-cystic growth pattern | 24
no vascular invasion | 24
renal capsule and adrenal gland were spared | 24
sarcomatoid differentiation | 24
large overlapping bundles of spindle-shaped cells | 24
tumor cells were negative for CD117 | 24
tumor cells were negative for CD10 | 24
tumor cells were negative for racemase | 24
tumor cells were negative for vimentin | 24
septic shock couldn't be controlled | 48
patient state deteriorated | 48
died | 72
chromophobe renal cell carcinoma | -672
abdominal pain | -672
hematuria | -672
abdominal mass syndrome | -672
decreased renal function | -672
proteinuria | -672
metastasis related pain | -672