29 years old | 0
female | 0
pregnant | 0
fever | -144
chills | -144
nonproductive cough | -144
breathlessness | -24
high-grade temperature | -144
rigor | -144
running nose | -144
sore throat | -144
postnasal drip | -144
malaise | -144
body ache | -144
lethargy | -144
weakness | -144
tachycardia | 0
tachypnea | 0
hypertension | 0
hypoxemia | 0
bilateral crackles | 0
bilateral nonhomogeneous opacity | 0
admitted to respiratory ICU | 0
H1N1 infection | 0
oseltamivir | 0
azithromycin | 0
paracetamol | 0
steroid prophylaxis | 0
fetal lung maturity | 0
transnasal humidified rapid-insufflation ventilatory exchange therapy | 0
high-risk consent | 0
surgery | 48
spinal anesthesia | 48
bupivacaine | 48
live birth | 48
uterotonics | 48
bilateral transversus abdominis plane block | 48
postoperative pain relief | 48
breathlessness | 48
noninvasive ventilator | 48
furosemide | 48
intensive care unit | 48
improved | 72
weaned off noninvasive ventilator | 72
discharged | 120