27 years old | 0
male | 0
fever | -48
presented to the clinic | 0
axillary temperature 101.8°F | 0
blood pressure 124/80 mmHg | 0
pulse 86 bpm | 0
denied prior comorbidities | 0
review of systems normal | 0
dengue NS1 test positive | 0
IgG/IgM negative | 0
haemoglobin 16.7 gm/dl | 0
white blood cell 6×10³/mm³ | 0
platelet 131×10³/mm³ | 0
unremarkable blood and urine investigations | 0
sent home with antipyretics | 0
two episodes of vomiting | 24
severe headache | 24
myalgia | 24
rash | 24
presented to the emergency room | 24
unwell appearance | 24
axillary temperature 100.5°F | 24
blood pressure 130/84 mmHg | 24
pulse 92 bpm | 24
petechiae over extremities, torso, abdomen, face | 24
platelet count trending down | 24
WBC count trending down | 24
mild hyponatremia (sodium 130 mEq/l) | 24
mild transaminitis | 24
hospitalized | 24
treated with analgesics | 24
treated with antipyretics | 24
treated with bed rest | 24
treated with fluids | 24
treated with nutritional support | 24
WBC dropped to 1900/mm³ | 144
platelet dropped to 48000/mm³ | 144
developed sharp chest pain | 144
chest pain aggravated during inspiration | 144
electrocardiogram normal | 144
Troponin-I normal | 144
ultrasonography revealed borderline splenomegaly | 168
ultrasonography revealed minimal left pleural effusion | 168
severe pain in lower limbs | 168
fever peaked at 100.4°F | 168
blood pressure 100/80 mmHg | 168
heart rate 97 bpm | 168
fever persisted | 168
pain became severe | 168
confined to bed | 168
focal tenderness in left buttock | 168
focal tenderness in left lumbosacral region | 168
focal tenderness in bilateral medial thigh | 168
no skin changes | 168
routine urine and stool examination normal | 168
urine culture no growth | 168
stool culture no growth | 168
blood culture no growth | 168
HIV negative | 168
Brucella negative | 168
Scrub Typhus negative | 168
Typhoid negative | 168
Malaria negative | 168
Leptospirosis negative | 168
NS1 test still positive | 168
IgG/IgM positive | 168
raised erythrocytic sedimentation rate (60 mm/h) | 168
raised C-reactive protein (90 mg/l) | 168
procalcitonin 0.29 ng/ml | 168
creatinine kinase normal | 168
troponin level normal | 168
echocardiography normal | 168
normal cannula site | 168
no recent trauma | 168
no intramuscular injections | 168
no recreational drug usage | 168
suspected intramuscular hematoma | 312
suspected secondary infection | 312
MRI ordered | 312
MRI showed left psoas muscle collection | 312
MRI showed left gluteal medius muscle collection | 312
MRI showed left adductor longus muscle collection | 312
MRI showed right pectineus muscle collection | 312
diffusion restriction within collections | 312
perilesional edema | 312
diagnosed pyomyositis | 312
started clindamycin | 312
started tazobactam-piperacillin | 312
upgraded to ICU | 312
aspirated purulent fluid from left adductor muscle | 312
gram staining negative | 312
culture grew Methicillin Sensitive Staphylococcus aureus | 312
sensitive to cloxacillin | 312
sensitive to tazobactam-piperacillin | 312
resistant to clindamycin | 312
acid fast bacilli stain negative | 312
PCR test for mycobacteria negative | 312
switched to cloxacillin | 312
switched to tazobactam-piperacillin | 312
received dual IV antibiotics for 2 weeks | 312
received oral cloxacillin for 4 weeks | 312
continuous clinical monitoring | 312
continuous USG monitoring | 312
repeat USG showed left adductor collection | 432
repeat USG showed left gluteal medius collection | 432
aspirated 30 ml pus-like fluid | 432
subsequent USG showed decreasing fluid | 432
discharged on oral antibiotics | 600
USG absence of intramuscular collection | 1008
