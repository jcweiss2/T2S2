48 years old | 0
    female | 0
    obesity | 0
    hypertension | 0
    referred for consideration of endoscopic sleeve gastroplasty | 0
    underwent endoscopic sleeve gastroplasty | 0
    general anesthesia | 0
    endoscopic suturing system | 0
    dual-channel endoscope | 0
    carbon dioxide insufflation | 0
    full thickness U-shaped suture pattern | 0
    placement of five sutures | 0
    immediate postoperative period | 0
    antiemetics | 0
    ondansetron | 0
    dimenhydrinate | 0
    dexamethasone | 0
    scopolamine | 0
    dipyrone | 0
    omeprazole | 0
    discharged | 24
    postoperative day 3 | 72
    abdominal pain | 72
    worsening abdominal pain | 96
    emergency department referral | 96
    fourth postoperative day | 96
    rigid abdomen | 96
    peritoneal irritation | 96
    leukocytosis | 96
    increased C-reactive protein | 96
    computed tomography free fluid in peritoneal cavity | 96
    biliary ascites | 96
    gallbladder puncture | 96
    emergent diagnostic laparoscopy | 96
    tubular stomach shape | 96
    peritoneal cavity lavage | 96
    gallbladder transfixed to stomach | 96
    biliary fluid collections | 96
    suture cut | 96
    laparoscopic cholecystectomy | 96
    intraoperative endoscopy | 96
    methylene blue test | 96
    intensive care unit admission | 96
    IV antibiotics | 96
    septic shock | 96
    discharge | 480
    weight loss | 4320
    no complications related to procedure | 4320
    