58 years old | 0
female | 0
hypertension | 0
admitted to the hospital | 0
fever | -120
dizziness | -120
denied dyspnea | -120
denied cough | -120
denied chills | -120
denied night sweats | -120
denied headache | -120
denied gastrointestinal symptoms | -120
no history of anorexia | 0
no history of weight loss | 0
born in the Dominican Republic | -175200
moved to New York City | -175200
denied use of tobacco | 0
denied use of alcohol | 0
denied use of recreational drugs | 0
febrile 39.5°C | 0
hypotensive | 0
blood pressure 88/40 mm Hg | 0
small cervical lymph nodes | 0
non-tender cervical lymph nodes | 0
soft cervical lymph nodes | 0
minimal bilateral rhonchi | 0
unremarkable abdominal exam | 0
unremarkable neurological exam | 0
unremarkable cardiac exam | 0
no organomegaly | 0
intact skin | 0
chest radiograph bilateral infiltrates | 0
admitted to intensive care unit | 0
severe sepsis | 0
pneumonia | 0
leukopenia 3.2 K/uL | 0
thrombocytopenia 144 K/uL | 0
elevated serum lactate dehydrogenase 1142 U/L | 0
IV ceftriaxone | 0
IV azithromycin | 0
persistent fever | 0
negative blood cultures | 0
negative urine cultures | 0
negative respiratory cultures | 0
negative AFB stains | 0
IV piperacillin-tazobactam | 0
IV vancomycin | 0
normal transthoracic echocardiogram | 0
CT chest bilateral infiltrates | 0
mediastinal lymphadenopathy | 0
subcarinal lymphadenopathy | 0
mild splenomegaly | 0
flexible fiber optic bronchoscopy | 144
bronchoalveolar lavage | 144
transbronchial biopsies | 144
EBUS-TBNA | 144
day 6 | 144
negative aerobic cultures | 144
negative AFB cultures | 144
negative fungal cultures | 144
negative viral cultures | 144
T cell lymphoma diagnosis | 144
CD4 positive | 144
CD3 positive | 144
CD43 positive | 144
BCL-2 positive | 144
CD20 negative | 144
CD10 negative | 144
CD79a negative | 144
PAX5 negative | 144
hypoxic respiratory failure | 360
intubation | 360
mechanical ventilation | 360
day 15 | 360
cervical lymph node excisional biopsy | 360
worsening cervical lymphadenopathy | 360
persistent fever | 360
peripheral T-cell lymphoma NOS | 360
CD3 positive | 360
CD4 positive | 360
CD5 positive | 360
CD43 positive | 360
Ki67 >90 positive | 360
CD20 negative | 360
CD79A negative | 360
CD7 negative | 360
CD15 negative | 360
bone marrow biopsy | 360
pancytopenia | 360
hemophagocytic lymphocytic histiocytosis | 360
negative AFB stains bone marrow | 360
negative fungal stains bone marrow | 360
tumor lysis syndrome | 360
acute renal failure | 360
hemodialysis | 360
rasburicase | 360
cyclophosphamide | 456
vincristine | 456
day 19 | 456
deterioration | 480
died | 480
day 20 | 480
AFB cultures cervical lymph nodes positive | 480
Mycobacterium tuberculosis complex | 480
AFB stains positive | 480
postmortem results | 480
