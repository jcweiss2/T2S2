46 years old | 0 | 0 
Asian-Indian | 0 | 0 
male | 0 | 0 
admitted to the hospital | 0 | 0 
tropical chronic pancreatitis | -8760 | 0 
oral pancreatic enzyme therapy | -8760 | 0 
non-insulin-dependent diabetes mellitus | -2190 | 0 
glucotrol | -2190 | 0 
midepigastric pain | -6 | 0 
pain control with narcotics | -6 | 0 
discharged | -48 | -48 
epigastric pain | 0 | 0 
nausea | 0 | 0 
vomiting | 0 | 0 
CT scan | 0 | 0 
fatty atrophy of pancreatic head and uncinate process | 0 | 0 
pancreatic duct filled with large calcifications | 0 | 0 
obstruction at the level of the neck | 0 | 0 
marked upstream ductal dilatation | 0 | 0 
admitted for management of pain | 0 | 0 
CT scan of the abdomen | -144 | -144 
chronic atrophic calcific pancreatitis | -144 | -144 
dilated pancreatic duct | -144 | -144 
intraductal calculi | -144 | -144 
ERCP | -144 | -144 
pancreatography | -144 | -144 
medically managed | -144 | -144 
discharged | -144 | -144 
fever | 48 | 48 
chills | 48 | 48 
rigors | 48 | 48 
severe sepsis | 48 | 48 
septic shock | 48 | 48 
transferred to the medical intensive care unit | 48 | 48 
intubated | 48 | 48 
hypoxemic respiratory failure | 48 | 48 
acute respiratory distress syndrome | 48 | 48 
multiorgan failure | 48 | 48 
broad-spectrum antibiotics | 48 | 240 
vasopressor support | 48 | 240 
activated recombinant human protein C | 48 | 240 
ultrasound of the abdomen | 48 | 48 
dilated pancreatic duct | 48 | 48 
calculus within the duct | 48 | 48 
diffusely echogenic pancreas | 48 | 48 
prominent common bile duct | 48 | 48 
bedside emergency ERCP | 72 | 72 
frank pus expelling spontaneously | 72 | 72 
evacuation of pus | 72 | 72 
cholangiogram | 72 | 72 
normal biliary tree | 72 | 72 
pancreatogram | 72 | 72 
marked dilatation of the main pancreatic duct | 72 | 72 
distal calculus | 72 | 72 
guide wire introduced | 72 | 72 
evacuation of pus | 72 | 72 
5-cm-long 5 F stent placed | 72 | 72 
reevaluation of the pancreas | 96 | 96 
contrast enhanced CT scan | 96 | 96 
inflammatory changes | 96 | 96 
edema | 96 | 96 
diminished dilatation of the pancreatic duct | 96 | 96 
distal migration of calculus | 96 | 96 
bilateral moderate pleural effusions | 96 | 96 
clinical improvement | 96 | 240 
stabilization of hemodynamic parameters | 96 | 240 
blood cultures grew Klebsiella ornithinolytica | 96 | 240 
extubated | 240 | 240 
transferred from the intensive care unit | 240 | 240 
completed antibiotic course | 240 | 240 
discharged home | 240 | 240 
follow-up examinations | 720 | 2160 
no further complications | 720 | 2160