58 years old | 0
female | 0
newly diagnosed AJCC stage IV metastatic melanoma | 0
metastatic spread to the lungs | 0
started on combination therapy nivolumab and ipilimumab | -432
received first two doses of nivolumab and ipilimumab | -432
arrived at emergency room | 0
severely altered | 0
hypotensive (66/41 mm Hg) | 0
tachycardic | 0
febrile (40.1 C) | 0
hypoxic (84% on room air) | 0
placed on BiPAP | 0
admitted to intensive care unit | 0
peripheral edema +3 in lower extremities extending to hips | 0
no significant past medical history | 0
elevated serum creatinine (2.8 mg/dL) | 0
elevated alanine transaminase (180 Units/L) | 0
elevated aspartate transaminase (165 Units/L) | 0
elevated lactate (10.9 mmol/L) | 0
elevated CRP (20.2 mg/L) | 0
mild leukocytosis (13.7 k/cumm) |-
chest X-ray showed pulmonary edema | 0
suspected septic shock | 0
met systemic inflammatory response syndrome criteria | 0
started on piperacillin-tazobactam | 0
started on vancomycin | 0
required norepinephrine | 0
required epinephrine | 24
required vasopressin | 24
continued BiPAP | 0
received fluids | 0
no improvement within 24 hours | 24
started on methylprednisolone | 24
concern for immune-mediated symptomology | 24
oxygenation saturation not maintained on BiPAP | 24
intubated | 24
no improvement after 2 days of methylprednisolone | 72
started on tocilizumab | 72
suspicion of CRS | 72
IL-6 levels measured | 72
TNF-α levels measured | 72
IL-6 level 21.4 pg/dL | 72
TNF1-α level 1,876 pg/dL | 72
oncology consulted | 72
tocilizumab chosen for CRS management | 72
consent obtained from family | 72
received 4 doses of tocilizumab | 72
received concurrent methylprednisolone | 72
symptoms did not improve | 72
trial of etanercept | 72
administration of etanercept | 72
symptoms improved | 72
extubated after 3 days | 168
improvement in laboratory results | 168
improvement in mental status | 168
improvement in fever | 168
discharged from hospital | 168
close follow-up with primary care provider and oncologist | 168
diagnosis of CRS stage 4 | 24
cytokine release syndrome | 24
fever | 0
hypotension | 0
hypoxia | 0
acute systemic inflammatory response | 0
multiple organ dysfunction | 0
activated T cells | 0
elevated interferon-gamma | 0
elevated IL-6 | 0
elevated TNF-α | 0
elevated IL-10 | 0
elevated IL-1 | 0
elevated IL-5 | 0
elevated IL-8 | 0
elevated macrophage colony-stimulating factors | 0
chills | 0
watery diarrhea | 0
activation of coagulation cascade | 0
vascular leakage | 0
lung injury | 0
cardiomyopathy | 0
activation of acute-phase proteins | 0
infection ruled out | 0
blood cultures | 0
empiric antibiotic therapy | 0
clinical diagnosis of CRS | 0
elevated CRP | 0
elevated ferritin | 0
elevated cytokine levels | 0
fever ≥38.0 C | 0
endo-organ dysfunction | 0
grade 4 CRS | 24
required vasopressors | 24
required intubation | 24
management with glucocorticoids | 24
management with tocilizumab | 72
management with etanercept | 72
refractory CRS | 72
tailored management based on cytokine levels | 72
elevated TNF-α | 72
trial of anakinra | 0
trial of siltuximab | 0
trial of ruxolitinib | 0
trial of baricitinib | 0
onset of CRS at first dose of immunotherapy | -432
awareness of CRS in clinicians | 0
patient education on CRS symptoms | 0
potential misdiagnosis as sepsis | 0
importance of measuring IL-6 and TNF-α | 72
need for guidelines in monoclonal antibody-induced CRS | 0
research on CRS treatment | 0
development of management guidelines | 0
written informed consent obtained | 0
no ethical approval required | 0
no conflicts of interest | 0
no funding required | 0
data availability statement | 0
mild leukocytosis (13.7 k/cumm) | 0
TNF-α level 1,876 pg/dL | 72
