81 years old | 0
male | 0
Caucasian | 0
admitted to the hospital | 0
fever | -504
progressive dyspnea | -504
dry cough | -504
left pleuritic chest pain | -504
chronic lymphocytic leukemia | -4018
Fludarabine treatment | -4018
Cyclophosphamide treatment | -4018
Rituximab treatment | -4018
type 2 diabetes mellitus | 0
hypertension | 0
hyperlipidemia | 0
chronic kidney failure | 0
eGFR of 28 mL/min/1.73 m2 | 0
no smoking | 0
no alcohol abuse | 0
worked as an upholsterer | 0
physical examination | 0
fever (38.1°C) | 0
tachycardia (105 bpm) | 0
peripheral percutaneous oxygen saturation was 100% | 0
tachypnea | 0
normal blood pressure | 0
almost abolished left vesicular murmur | 0
no adenopathy | 0
no hepatomegaly | 0
no splenomegaly | 0
normal cardiovascular examination | 0
normal neurologic examination | 0
neutrophilia (18.7 g/L) | 0
elevated CRP (297 mg/L) | 0
stable lymphocytosis (242 g/L) | 0
anemia (7.8 g/L) | 0
large left pleural effusion | 0
contralateral tracheal deviation | 0
walled-off, loculated left pleural effusion | 0
normal right lung parenchyma | 0
citrine exudate | 0
pleural protein 37 g/L | 0
pleural fluid protein to serum ratio 0.61 | 0
intravenous treatment with cefotaxime | 0
persistence of fever | 24
persistence of neutrophilia | 24
severe hypoxemia | 24
bacteriological standard culture of the pleural liquid sample was negative | 24
repeated blood cultures were negative | 24
auramine stained sputum smears and cultures were negative | 24
spot-test for tuberculosis was not performed | 0
surgical thoracentesis | 240
evacuation of 2 liters of purulent liquid | 240
thick and nodular pleura | 240
white pseudo-membranes | 240
treatment with metronidazole | 240
cytobacteriological examination and cultures of the liquid were negative | 240
lymphocyte phenotyping ruled out B-cell lymphoma | 240
multiple organ failure | 264
intensive care unit admission | 264
antibiotherapy with cefepime and amikacin | 264
invasive mechanical ventilation | 264
vasopressor infusion | 264
renal replacement therapy | 264
uncontrolled septic shock | 264
death | 288
mycobacterial culture of surgical pleural samples yielded Gram-negative bacilli | 288
L. pneumophila identified | 288
L. pneumophila serogroup 1 | 288
urinary antigen research confirmed the presence of L. pneumophila serogroup 1 | 288
male sex | 0
aged more than 50 years | 0
chronic lymphocytic leukemia with history of immunocompromising treatments | 0
chronic kidney failure | 0
diabetes mellitus | 0
weaned smoking | 0
pleural empyema | 0
L. pneumophila infection | 0
sepsis | 0
septic shock | 264
multiple organ failure | 264
uncontrolled sepsis | 288
L. pneumophila serogroup 1 pleural empyema | 288