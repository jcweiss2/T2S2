47 years old | 0
female | 0
poorly controlled type 1 diabetes mellitus | -672
heart failure | -672
mild severe acute coronavirus respiratory virus-2 | -1344
left lower extremity deep vein thrombosis | -672
altered mental status | 0
burning sensation of her left hand | 0
cachectic | 0
alert to self | 0
comfortable | 0
blood pressure of 104/65 mm/Hg | 0
pulse of 88 beats/min | 0
respiratory rate of 20 breaths/min | 0
oxygen saturation of 99% on room air | 0
wet gangrene of the left fourth digit | 0
leukocytosis | 0
acute kidney injury | 0
diabetic ketoacidosis | 0
glucose of 746 mg/dl | 0
anion gap of 30 | 0
atrophy of the fourth digit with subcutaneous gas | 0
consolidative and reticular opacities in the right lower lung | 0
cavitary right lower lobe lesion with possible reversed halo sign | 0
vancomycin | 0
piperacillin-tazobactam | 0
clindamycin | 0
admitted to the intensive care unit | 0
resolution of DKA | 48
amputation of her left fourth digit | 48
left wrist disarticulation | 48
worsening leukocytosis | 72
white blood cell count of 54,320 | 72
broadened antimicrobial coverage | 72
vancomycin | 72
meropenem | 72
doxycycline | 72
liposomal amphotericin B | 72
bronchoscopy | 72
infiltrates of the right middle and lower lobe | 72
diffuse necrotic tissue | 72
fibrinous clot | 72
thoracic surgery | 72
operative management | 72
right lower lobectomy | 96
posaconazole | 96
bilateral frontal lobe punctate infarcts | 96
right atrial vegetation | 96
patent foramen ovale | 96
AngioVac extraction | 120
small vegetation | 120
no tissue obtained for culture or pathology | 120
bronchoalveolar lavage cytologic specimen | 168
pauciseptate hyphae of a zygomycete | 168
Rhizopus species | 168
hand surgical pathology | 168
hyphae present within vessels and around nerves | 168
vascular spread | 168
cutaneous inoculation | 168
stable post-operatively | 168
transferred to the general medicine floor | 168
re-admitted to the ICU | 240
hypothermia | 240
hypotension | 240
vasopressor support | 240
acute metabolic encephalopathy | 240
bilateral pleural effusions | 240
percutaneous drains | 240
acute kidney injury | 240
mixed transaminitis | 240
antifungal medications | 240
discontinue further treatment | 336
comfort care | 336
passed away | 360