56 years old | 0
    male | 0
    admitted to the hospital | 0
    scrotal pain | -96
    myalgia | -96
    inability to walk | -96
    alcohol abuse | 0
    40 pack-year smoking history | 0
    fulminant necrosis of the scrotum | 0
    necrosis of the dorsum of both feet | 0
    necrosis of the heels of both feet | 0
    necrosis of the left middle finger | 0
    intravenous benzylpenicillin | 0
    flucloxacillin | 0
    transferred to the nearest regional center | 0
    diagnosis of scrotal Fournier gangrene | 0
    concurrent multifocal necrotizing fasciitis | 0
    intravenous clindamycin | 0
    meropenem | 0
    vancomycin | 0
    surgical exploration | 0
    debridement | 0
    global necrosis of scrotum | 0
    copious purulent discharge | 0
    bilateral nonviable testes | 0
    scrotal debridement | 0
    bilateral orchiectomy | 0
    debridement of necrotic tissue from both feet | 0
    debridement of necrotic tissue from left middle finger | 0
    admitted to the intensive care unit | 0
    intubated | 0
    intravenous vasopressor support (noradrenaline) | 0
    antibiotics | 0
    scrotal tissue culture revealed Streptococcus intermedius | 0
    scrotal tissue culture revealed Escherichia coli | 0
    scrotal tissue culture revealed Klebsiella oxytoca | 0
    scrotal tissue culture revealed Staphylococcus aureus | 0
    histological examination of limb tissue consistent with necrotizing fasciitis | 0
    spent 6 days in ICU | 24
    spent 4 days on noradrenaline vasopressor support | 24
    spent 24 days on the surgical ward | 24
    scrotal debridement on day 2 | 48
    left medial thigh exploration on day 2 | 48
    insertion of bilateral middle ear ventilation tubes on day 2 | 48
    scrotal wound reexploration and closure on day 8 | 192
    further debridement of limb wounds on day 8 | 192
    further debridement on day 16 | 384
    split skin grafts from the left thigh to bilateral heel wounds on day 16 | 384
    use of vasopressors | 0
    discharged on day 30 | 720
    scrotal wound stabilized | 720
    bilateral skin grafts showed good uptake | 720
    oral ciprofloxacin | 720
    amoxicillin/clavulanate | 720
    lifelong testosterone replacement therapy | 720
    discharged home after 60 days of inpatient rehabilitation | 1440
    full recovery | 1440
    well 5 months on from initial presentation | 3600
    plans to return to fruit picking | 3600
    