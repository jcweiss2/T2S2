67 years old | 0
male | 0
admitted to the hospital | 0
history of worsening dyspnea | -96
irritating cough | -96
expectoration of brownish sputum | -96
general weakness | -96
metabolic syndrome | 0
diabetes | 0
hyperlipidemia | 0
PPI | 0
subfebrile | 0
nausea | 0
no vomiting | 0
no diarrhea | 0
no chest pain | 0
no loss of taste | 0
no loss of smell | 0
blood saturation 92% O2 | 0
borderline blood pressure 115/60 mm Hg | 0
mild tachycardia 100 rpm | 0
rapid test for COVID-19 positive | 0
PCR test for COVID-19 positive | 0
bilateral pneumonia | 0
elevation of inflammatory markers | 0
decompensated diabetes mellitus | 0
normal renal function | 0
normal liver function | 0
antibiotic therapy | 0
corticoids | 0
bronchodilators | 0
LMWH | 0
adjustment of diabetic medication | 0
shortness of breath | 24
irritating cough | 24
desaturation up to 76% O2 | 24
transfer to intensive care unit | 24
HFNO therapy | 24
continuation of corticoids and antibiotics | 24
increase of LMWH dose | 24
severe hypoxemia | 144
arterial astrup blood gas analysis | 144
indication for translation to anesthesiology and resuscitation department | 144
intubation | 144
construction of tracheostomy | 144
escalation of ATB | 144
nutrition via nasogastric tube | 144
circulatory support of vasopressors | 144
septic shock | 144
withdrawal of catecholamines | 240
subsidence of febrile episodes | 240
decrease of inflammatory markers | 240
discontinuation of sedatives | 240
regain of consciousness | 240
low muscle strength | 240
considered noninfectious | 504
planned transfer to rehabilitation care ward | 504
sudden rapid deterioration | 552
circulatory instability | 552
tachypnea | 552
fibrillation | 552
massive enterorrhagia | 552
drop of hemoglobin to 81 g/L | 552
septic shock | 552
intubation | 552
circulatory resuscitation | 552
administration of catecholamines | 552
multiple blood substitutes | 552
hemostatic therapy | 552
discontinuation of LMWH therapy | 552
abdominal ultrasound | 552
undilated small-bowel loops | 552
meteoric colon | 552
no obvious wall thickening | 552
no free fluid in abdominal cavity | 552
gastrofibroscopy | 552
colonoscopy | 552
normal mucosa from esophagus to D2 part of duodenum | 552
no signs of bleeding | 552
clarity of colon wall aggravated | 552
presence of intestinal contents and coagula | 552
no source of bleeding or mural lesion | 552
CT angiography of abdomen | 552
liquid content in cecum | 552
suspected coagulum in sigmoid colon and ampulla recti | 552
distended cecum and sigmoideum | 552
no wall thickening | 552
no clear source of bleeding | 552
indication for acute abdominal revision | 552
midline laparotomy | 552
distended colon | 552
translucent hemorrhagic filling | 552
desufflation of cecum | 552
revision of small intestine | 552
enterotomy in terminal ileum | 552
no signs of bleeding | 552
right-sided hemicolectomy | 552
ileotransversoanastomosis | 552
histological examination | 552
ischemic enteritis and colitis | 552
mucosal ulcerations | 552
no infectious or IBD inflammation | 552
no Dieulafoy lesion | 552
no dysplasia or malignancy | 552
stabilization of patient's condition | 624
weaning | 624
adjustment of intestinal passage | 624
enteral nutrition via nasogastric probe | 624
transfer to post-acute intensive care unit | 1008
readmission for recurrent GIT bleeding | 1344
colonoscopy | 1344
small ulceration in area of ileotransversoanastomosis | 1344
conservative management with hemodynamic therapy | 1344
transfer back to post-acute intensive care department | 1344