46 years old | 0
male | 0
ulcerative colitis | -72
malaise | -72
fever | -72
loss of appetite | -72
presented to emergency department | 0
blood pressure 124/46 mmHg | 0
heart rate 122 beats per min | 0
SpO2 98% | 0
respiratory rate 16/min | 0
body temperature 40.2°C | 0
alert | 0
lying in bed | 0
chills | 0
nausea | 0
cardiac arrest | 0
chest compression | 0
tracheal intubation | 0
ECG ventricular fibrillation | 0
defibrillation | 0
adrenaline administered | 0
resuscitated | 0
diagnosed Brugada syndrome | 0
ECG coved-type ST elevation V1 V2 | 0
fever subsided with acetaminophen | 24
hypercalcemia 14.8 mg/dL | 0
admitted to intensive care unit | 0
hypotension | 0
suspected septic shock | 0
CT high-density area descending colon | 0
increased lactate level | 0
increased white blood cell count | 0
increased procalcitonin level | 0
initiated tazobactam-piperacillin | 0
initiated vasopressors | 0
extubation | 48
fever recurrence | 120
contrast-enhanced CT liver abscess | 120
changed antibiotics to meropenem | 120
changed antibiotics to vancomycin | 120
maintained antibiotics for 3 weeks | 120
performed puncture drainage | 120
infection controlled | 720
positive pilsicainide test | 720
ICD implantation | 720
discharged | 720
family history sudden death | 0
hypercalcemia causes examined | 0
high parathyroid hormone levels | 0
Tc scintigraphy anterior mediastinum uptake | 0
tumor resection post-discharge | 720
followed up ECG | 720
followed up serum calcium | 720
ectopic parathyroid adenoma | 720
CT pituitary tumors | 720
MRI adrenal tumors | 720
nonfunctional pituitary adenomas | 720
nonfunctional adrenal tumors | 720
diagnosed multiple endocrine neoplasia type 1 | 720
consent obtained | 0
