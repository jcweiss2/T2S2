57 years old | 0
female | 0
hypertension | -672
recurrent cystitis | -672
type 2 diabetes mellitus | -672
ESRD | -672
hemodialysis | -672
lethargic | -12
barely conscious | -12
fever | -12
temperature of 95.5F | 0
heart rate 102 beats per minute | 0
respiratory rate 10 cycles per minute | 0
blood pressure 76/55 mmHg | 0
soft abdomen with mild distension | 0
trace pedal edema | 0
intubated | 0
admitted to MICU | 0
leukocytosis | 0
normocytic anemia | 0
lactic acidosis | 0
elevated serum creatinine levels | 0
hemoglobin A1C level 6.1% | 0
arterial blood gas levels normal | 0
urinalysis positive for bacteria | 0
urinalysis positive for leukocyte esterase | 0
urinalysis positive for nitrites | 0
abdominopelvic CT scan showed extensive small and large bowel thickening | 0
abdominopelvic CT scan showed thickening and irregularity of the bladder wall | 0
abdominopelvic CT scan showed mild ascites | 0
chest X-ray normal | 0
brain CT scan normal | 0
initiated on IV fluids | 0
initiated on empiric IV antibiotics | 0
initiated on norepinephrine | 0
initiated on continuous renal replacement therapy | 0
general surgery team consulted | 0
evaluated for possible complicated ischemic colitis | 0
presumptive diagnosis of ischemic colitis with bacteremia | 0
no acute surgical intervention warranted | 0
clinical condition deteriorated | 24
persistently febrile | 24
tachycardic | 24
requiring more doses of norepinephrine | 24
abdomen more distended | 24
laboratory parameters worsened | 24
blood microbiology studies resulted for Escherichia coli | 24
urine microbiology studies resulted for Escherichia coli | 24
taken to operating room for urgent exploratory laparotomy | 24
suspected peritonitis from colon ischemia | 24
laparotomy revealed necrotic and ruptured bladder wall | 24
free fluid in abdominopelvic cavity | 24
no bowel ischemia or perforation | 24
partial cystectomy | 24
pathologic analysis confirmed bladder tissue inflammation and necrosis | 24
no malignancy | 24
withdraw life support treatment and care | 96
died | 107