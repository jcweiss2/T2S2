88 years old | 0
    male | 0
    presented to the emergency room | 0
    skin color change in the right scrotal area | -24
    right scrotal pain | -168
    right scrotal swelling | -168
    administered oral fluoroquinolone | -168
    administered ciprofloxacin | -168
    symptoms aggravated | -168
    skin color changed from red to black | -24
    foul-smelling | -24
    visited the urology department for voiding dysfunction | -62760
    a-blocker (silodosin 8 mg daily) | -62760
    5 alpha reductase inhibitor (finasteride once daily) | -62760
    voiding symptom aggravated | -62760
    total IPSS score 26 | -62760
    Quality of Life score 5 | -62760
    maximal flow rate (Qmax) 6.5 mL/sec | -62760
    voiding volume 182 mL | -62760
    residual urine volume 258 mL | -62760
    prostate volume 126 cc | -62760
    diagnosed with refractory to medical therapy | -62760
    planned TURP | -62760
    not suited for surgery under general anesthesia | -62760
    high ASA score (grade III) | -62760
    history of NSTEMI | -62760
    cerebrovascular accident | -62760
    poor-controlled COPD | -62760
    spinal anesthesia contraindicated due to spinal stenosis | -62760
    decided MIS under local anesthesia | -62760
    intraurethral lidocaine injection | -62760
    analgesic injection intravenously | -62760
    implanted Memokath 028 | -62760
    Qmax 14.8 mL/sec after 6 months | -57600
    residual urine volume 85 mL after 6 months | -57600
    suprapubic cystostomy | -35040
    prostatic stent not working | -35040
    blood pressure 110/70 mmHg | 0
    heart rate 90/min | 0
    body temperature 36.0°C | 0
    oxygen saturation 96% | 0
    skin necrosis right lower abdomen to right scrotum | 0
    left lower abdomen normal | 0
    left scrotum normal | 0
    penis normal | 0
    digital rectal examination tenderness | 0
    digital rectal examination heat of entire prostate | 0
    elevated white blood cell count 13.62 /uL | 0
    elevated C-reactive protein 23.79 mg/dL | 0
    elevated procalcitonin 7.12 ng/mL | 0
    elevated serum lactate 3.5 mmol/L | 0
    elevated serum creatinine 2.47 mg/dL | 0
    elevated serum glucose 133 mg/dL | 0
    pyuria | 0
    Enterobacter cloacae isolated in urine | 0
    Enterobacter cloacae isolated in blood | 0
    Fournier’s gangrene severity index 7 points | 0
    serum potassium 5.5 | 0
    serum creatinine 2.47 | 0
    serum bicarbonate 16.3 | 0
    emphysematous changes on CT | 0
    inflammatory infiltration on CT | 0
    prostatic urethral stent observed | 0
    enlarged prostate | 0
    no abscess formation | 0
    no emphysematous change in prostate and urethra | 0
    Fournier’s gangrene | 0
    acute prostatitis | 0
    started meropenem | 0
    started vancomycin | 0
    started clindamycin | 0
    necrotic tissues excised | 0
    right orchiectomy performed | 0
    necrotic change of right spermatic cord | 0
    necrotic change of epididymis | 0
    culture swab in open wound | 0
    Memokath 028 stent removed | 0
    erythematous change of prostatic urethra | 0
    vital sign unstable | 0
    persisted low blood pressure | 0
    tachycardia | 0
    admitted to ICU | 0
    mechanical ventilation | 0
    broad-spectrum antibiotics continued | 0
    total parenteral nutrition | 0
    hemodialysis initiated | 24
    incomplete surgical debridement | 0
    necrotic tissues debrided several times | 0
    follow-up culture negative | 0
    elevated liver enzyme | 288
    elevated bilirubin | 288
    decreased platelet count 23000/L | 312
    prolonged prothrombin time | 312
    prolonged international normalized ratio | 312
    died | 336
    multiorgan failure | 336
    sepsis | 336