63 years old | 0
woman | 0
admitted to the ICU | 0
alcohol use disorder | 0
type 2 diabetes mellitus | 0
hypertension |.0
chronic pancreatitis | 0
pseudocyst | 0
mixed hemorrhagic/distributive shock | 0
acute gastrointestinal bleed | 0
diabetic ketoacidosis | 0
lethargic | -24
declining responsiveness | -24
hypothermic to 32.4°C | -24
hypotensive with blood pressure 52/33 mmHg | -24
hemoglobin 13 g/dL | -24
glucose >1500 mg/dL | -24
beta-hydroxybutyrate >22.50 mmol/L | -24
creatinine 3.55 mg/dL | -24
BUN 101 mg/dL | -24
bicarbonate 5 mmol/L | -24
pH 7.01 | -24
large-volume hematemesis | -24
requiring 2 units packed red blood cells | -24
intubation | -24
airway protection | -24
placement of right internal jugular vein central line | -24
started on insulin | -24
started on pantoprazole drips | -24
given 1 dose of 2g i.v. ceftriaxone | -24
transferred to our hospital | -24
afebrile | 0
tachycardic 120 bpm | 0
mean arterial pressure 90/60 mmHg | 0
norepinephrine infusion | 0
vasopressin infusion | 0
pH 7.21 | 0
bicarbonate 22 mmol/L | 0
glucose 902 mg/dL | 0
anion gap 28 mmol/L | 0
potassium 3.7 mmol/L | 0
BUN 84 mg/dL | 0
creatinine 2.47 mg/dL | 0
lipase 69 U/L | 0
C-reactive protein 262 mg/L | 0
sedimentation rate >120 mm/h | 0
undetectable ethanol | 0
hemoglobin 15 g/dL | 0
platelets 165000 per cu mm | 0
white blood cell count 3300 per cu mm | 0
infectious diseases workup | 0
blood cultures | 0
sputum cultures | 0
urine cultures | 0
chest X-ray showed bilateral lower lung patchy opacities | 0
remained on norepinephrine | 0
remained on vasopressin | 0
remained on insulin drips | 0
started on piperacillin/tazobactam | 0
blood cultures positive for Candida species | 24
started on micafungin | 24
cultures speciated to C. albicans | 24
blood cultures on days 1-3 | 24
blood cultures grew C. glabrata on days 5 and 7 | 120
line holiday | 24
removal of arterial line | 24
removal of right internal jugular vein central line | 24
transthoracic echocardiogram | 24
CT chest | 24
CT abdomen and pelvis | 24
ophthalmologic exam | 24
left hip hemiarthroplasty | 0
plain films | 24
attempted hip aspiration | 24
upper and lower extremity duplexes | 168
DVT in right internal jugular vein | 168
started on heparin drip | 168
clearance of clot | 240
clearance of blood cultures | 240
remained on fluconazole | 168
planned 3 months of enoxaparin | 168
stayed in hospital 31 days | 744
discharged to skilled nursing facility | 744
