53 years old | 0
male | 0
hypertension | 0
diabetes mellitus | 0
hypothyroidism | 0
stable dilated cardiomyopathy | 0
admitted to the hospital | 0
prolonged pyrexia | 0
coronary angiography | -1344
normal coronary anatomy | -1344
moderate- to high-grade fever | -1128
standard investigations | -1128
routine blood cultures | -1128
imaging | -1128
transferred to our care | -2016
febrile | -2016
toxic | -2016
early diastolic murmur in the aortic area | 0
hemoglobin 8.3 g/dL | 0
white blood cells 9200 cells/mm³ | 0
platelets 223000/mm³ | 0
serum creatinine level 2.2 mg/dL | 0
erythrocyte sedimentation rate 88 mm/h | 0
urine analysis showed 3-5 RBCs/hpf | 0
raised 24-h urine protein of 1527 mg/24 h | 0
ultrasonography kidney sizes normal | 0
no evidence of pyelonephritis or abscess | 0
mild hepatosplenomegaly | 0
no evidence of focal lesions in the spleen or liver | 0
chest roentgenogram mildly prominent pulmonary vasculature | 0
cardiomegaly | 0
no significant lung parenchymal pathology | 0
2D ECHO LVEF 30% | 0
normal heart valves | 0
global hypokinesia | 0
repeat 2D echo mild aortic regurgitation | 0
three discrete small mobile vegetations on aortic valve | 0
no evidence of cusp perforation or ring abscess | 0
other cardiac valves normal | 0
LVEF 20% | 0
transesophageal echo confirmed findings | 0
choroidal infiltrates | 0
no evidence of embolization to skin or other organs | 0
anti-ANA negative | 0
anti-dsDNA antibody negative | 0
anti&ndash;ANCA negative | 0
complement levels (C3 and C4) normal | 0
thyroid profile normal | 0
treated for heart failure | 0
started on ceftriaxone | 0
routine serial bacterial blood cultures | 0
BACTEC Myco/F Lytic medium demonstrated NTM | 0
linezolid added | 0
clarithromycin added | 0
species identification revealed M. abscessus | 0
drug sensitivities obtained | 0
sensitive to amikacin | 0
sensitive to clarithromycin | 0
sensitive to linezolid | 0
sensitive to tobramycin | 0
intermediate sensitivity to cefoxitin | 0
resistant to doxycycline | 0
resistant to imipenem | 0
resistant to cefepime | 0
resistant to ceftriaxone | 0
resistant to minocycline | 0
resistant to amox&ndash;clavulanic acid | 0
linezolid continued | 0
clarithromycin continued | 0
isoniazid added | 0
ethambutol added | 0
cefoxitin added | 0
defervesced after 7 weeks | 168
linezolid withheld | 168
bone marrow suppression | 168
linezolid reinstituted | 528
after 3 weeks therapy | 504
creatinine stabilized at 2.6 mg/dL | 504
previous peak creatinine 3.6 mg/dL | 504
dyspnea improved | 504
repeat 2D echo LVEF 40% | 504
valvular vegetations present | 504
blood cultures still grew mycobacteria | 504
aortic valve replacement surgery considered | 504
withheld due to comorbidities | 504
patient reluctance to undergo procedure | 504
repeat 2D ECHO at 4 weeks | 672
no change in vegetation size | 672
discharged on antimycobacterial antibiotics | 672
subsequently developed worsening cardiac failure | 672
died of pulmonary edema | 672
renal dysfunction | 672
hypothyroidism |*Annotation*
