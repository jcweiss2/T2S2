64 years old| 0
male| 0
admitted to the hospital| 0
COVID-19| 0
asymptomatic sinus bradycardia| 0
heart rate 30-45 BPM| 0
right heart axis| 0
incomplete right bundle branch block| 0
QRS 100, 120 msec| 0
downsloping depression of ST-segment| 0
T inversion| 0
normotensive| 0
blood pressure 135/54| 0
good pulse volume| 0
oxygen saturation 98-99%| 0
jugular venous pressure not raised| 0
no radio-radial delay| 0
no radio-femoral delay| 0
pansystolic murmur grade III| 0
moderate aortic regurgitation| 0
thickened aortic valve| 0
dilated left ventricular chamber| 0
ejection fraction 70%| 0
no pericardial effusion| 0
pulmonary artery systolic pressure 10.0+5.0 mmHg| 0
no foot oedema| 0
baseline haematological parameters within normal limits| 0
baseline biochemical parameters within normal limits| 0
intravenous atropine 0.5 mg| 0
unsuccessful| 0
intravenous dopamine 5 mg| 0
uptitrated to 15 mg| 0
no improvement in heart rate| 0
persistent wide pulse pressure| 0
transcutaneous cardiac pacing| 0
dopamine weaned off| 0
noradrenaline infusion titrated| 0
heart rate improved to 45-60 BPM| 24
systolic blood pressure 110-150 mmHg| 24
diastolic blood pressure 60-90 mmHg| 24
blood pressure decreased to 88/54 mmHg| 96
heart rate 54 BPM| 96
transvenous pacing via subclavian access| 96
heart rate setting 80| 96
output 10| 96
shortness of breath| 96
chest pain| 96
sweating| 96
pacer removed| 96
re-implantation via jugular access| 96
lower abdominal pain| 96
no bowel movements since admission| 96
vomited once| 96
streaks of blood on diapers| 96
severe metabolic acidosis| 96
pH 7.013| 96
pO2 71.9| 96
pCO2 43.5| 96
HCO3- 11.0| 96
anion gap 33.1 mEq/l| 96
free-flow gastric decompression 665 ml| 96
yellowish faecal material| 96
computed tomography abdomen| 96
short segment circumferential wall thickening| 96
proximal ascending colon| 96
inflammatory changes| 96
infective changes| 96
right inguinal hernia| 96
small bowel obstruction| 96
mesenteric content| 96
proximal bowel dilatation| 96
right inguinal hernia soft| 96
reducible| 96
non-tender| 96
measuring 7x5 cm| 96
no overlying skin changes| 96
no surgical intervention| 96
clinical condition deteriorated| 96
multiorgan failure| 96
persistent hyperglycaemia| 96
Dextrostix 14.0 mmol/l| 96
cardiorenal syndrome| 96
anuria| 96
worsening metabolic acidosis| 96
urea 16.5 mmol/l| 96
creatinine 343 µmol/l| 96
fulminant hepatic failure| 96
ALT 4,944 U/l| 96
AST 16,722 U/l| 96
hyperbilirubinemia| 96
total bilirubin 63 µmol/l| 96
thrombocytopaenia| 96
platelet count 73x103/µl| 96
coagulopathy| 96
NAC regimen| 96
third space loss| 96
global pericardial effusion| 96
2.0-2.5 cm| 96
right ventricular wall thickness| 96
double strengths of triple inotropic support| 96
haemodialysis| 96
SLEDD| 96
CVVH| 96
fresh-frozen plasma| 96
packed cells| 96
platelet concentrate| 96
empirical antibiotics escalated to meropenem| 96
succumbed to disease| 144
