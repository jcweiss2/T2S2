52 years old | 0 | 0 
male | 0 | 0 
body mass index of 23.6 kg/m2 | 0 | 0 
no comorbidities | 0 | 0 
admitted to the hospital | 0 | 0 
open modified Scopinaro procedure | -7440 | -7440 
weight of 216 kg | -7440 | -7440 
BMI 57.4 kg/m2 | -7440 | -7440 
weight reganance | -2400 | -1680 
incisional hernia | -2400 | -1680 
bariatric revisional surgery | -1680 | -1680 
hernia repair | -1680 | -1680 
gastric pouch leak | -1680 | -840 
multiple intra-abdominal collections | -1680 | -840 
sepsis | -1680 | -840 
conservative management | -1680 | -840 
open abdomen | -1680 | -840 
negative wound pressure therapy | -1680 | -840 
parenteral nutrition | -1680 | -840 
intravenous antibiotics | -1680 | -840 
epithelized gastrocutaneous fistula | -840 | 0 
controlled but persistent drainage | -840 | 0 
upper endoscopy | -24 | 0 
fistulous orifice | -24 | 0 
extraluminal extravasation | -24 | 0 
recurrent left subphrenic abscess | -24 | 0 
endoscopic treatment | 0 | 0 
argon plasma coagulation | -720 | -720 
internal and external drainages | -720 | -720 
clipping | -720 | -720 
fibrin sealants | -720 | -720 
e-vac therapy | -720 | -720 
stenting | -720 | -720 
multidisciplinary team discussion | 0 | 0 
decision to proceed with an innovative endoscopic technique | 0 | 0 
placement of a CSDO | 0 | 0 
Occlutech muscular VSD occluder | 0 | 0 
procedure performed in the catheterization laboratory | 0 | 2 
intravenous sedation | 0 | 2 
topic anesthesia | 0 | 2 
fistula cannulated | 0 | 2 
extraluminal leakage documented | 0 | 2 
Amplatz extra stiff guidewire | 0 | 2 
delivery system introduced | 0 | 2 
CSDO deployed | 0 | 2 
contrast study | 2 | 2 
no extravasation of contrast material | 2 | 2 
restricted oral intake | 2 | 26 
liquid diet | 26 | 240 
regular diet | 240 | 240 
pigtail drain positioned | 240 | 1008 
accidental displacement of the pigtail | 1008 | 1008 
systemic signs of sepsis | 1008 | 1008 
computed tomography | 1008 | 1008 
fluoroscopy | 1008 | 1008 
recurrence of the abscess | 1008 | 1008 
partial dislodgment of the 8-mm mVSD CSDO | 1008 | 1008 
second attempt with an oversized disc | 1008 | 1010 
Occlutech Figulla Flex II UNI 24-mm | 1010 | 1010 
sealing of the fistulous orifice | 1010 | 1010 
6-month clinical and imaging follow-up | 3024 | 3024 
upper endoscopy | 3024 | 3024 
contrast-enhanced CT scan | 3024 | 3024 
device engrafted | 3024 | 3024 
reduction of the chronic abscess | 3024 | 3024 
no signs of fistula recurrence | 3024 | 3024 
pigtail removed | 3024 | 3024 
no drainage observed | 3024 | 3024