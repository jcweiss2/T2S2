57 years old | 0
female | 0
admitted to the hospital | 0
acute abdominal pain | -72
abdominal pain aggravated after ingestion of food | -72
palpitation | -72
vomiting | -72
no stool or flatus | -48
chronic smoker | -8760
Chronic Obstructive Pulmonary Disease | -8760
medication for Chronic Obstructive Pulmonary Disease | -8760
tachycardia | 0
sinus rhythm | 0
oxygen saturation 85% | 0
blood pressure 95/70 mmHg | 0
body temperature 38.7°C | 0
respiratory rate 22 breaths/min | 0
COVID-19 positive | 0
leukocytosis | 0
raised amylase | 0
liver function test abnormal | 0
metabolic acidosis | 0
raised lactate level | 0
nasogastric tube decompression | 0
Foley catheterization | 0
crystalloids administered | 0
supplemental oxygen | 0
analgesics administered | 0
intravenous antibiotics | 0
emergency laparotomy | 12
gangrenous small bowel | 12
resection of gangrenous segment | 12
double barrel loop ileostomy | 12
Meropenem IV | 24
Vancomycin IV | 24
low molecular weight Heparin | 24
total parenteral nutrition | 24
COVID pneumonia | 144
reintubation | 144
sepsis | 168
Acute Kidney Injury | 168
multi-organ dysfunction syndrome | 168
expired | 336
D-dimer elevated | 0
fibrinogen elevated | 0
thromboembolism prophylaxis | 0 
anticoagulant use | 24 
histopathological report showed small bowel necrosis | 24 
microthrombi in the lamina propria | 24 
microthrombi in the submucosa | 24 
glandular necrosis | 24 
mucosal denudation | 24 
decreased crypts in the lamina propria | 24 
submucosa edematous | 24 
dense acute inflammatory cells | 24 
hyalinized blood vessels | 24 
microthrombi formation | 24 
abdominal X-ray showed prominent dilated small bowel loops | 0
abdominal X-ray showed multiple air fluid levels | 0
CECT scan showed collection of fluid | 0
CECT scan showed patent mesenteric vessels | 0 
non-occlusive mesenteric ischemia | 12 
acute mesenteric ischemia | 12 
small intestinal hypoperfusion | 12 
bowel wall necrosis | 12 
endothelial inflammation | 0
thrombin formation | 0
complement activation | 0
immune response initiation | 0 
vasopressors | 0
hemodynamic instability | 0
metabolic derangements | 0
positive pressure ventilation | 0
viral enteritis | 0 
percutaneous endovascular thrombectomy | 0 
thromboembolism | 0 
anticoagulation | 24 
in-hospital mortality risk | 0 
prognosis | 0 
mortality | 336 
informed consent | -72 
publication of case report | -72 
accompanying images | -72 
written consent | -72 
Editor-in-Chief | -72 
review | -72 
ethical approval | -72 
funding | -72 
grant | -72 
public sector | -72 
commercial sector | -72 
not-for-profit sector | -72 
guarantor | -72 
research registration | -72 
CRediT authorship | -72 
conceptualization | -72 
supervision | -72 
writing | -72 
original draft | -72 
review and editing | -72 
conflict of interest | -72 
acknowledgments | -72 
patient | -72 
colleagues | -72 
insightful comments | -72 
Muna Sharma | -72 
Subodh Dhakal | -72 
colleagues | -72 
insightful comments | -72 
patient | -72 
acknowledgments | -72 
conflict of interest | -72 
CRediT authorship | -72 
research registration | -72 
grant | -72 
funding | -72 
ethical approval | -72 
review | -72 
written consent | -72 
Editor-in-Chief | -72 
publication of case report | -72 
accompanying images | -72 
informed consent | -72 
prognosis | 0 
in-hospital mortality risk | 0 
anticoagulation | 24 
thromboembolism | 0 
percutaneous endovascular thrombectomy | 0 
viral enteritis | 0 
positive pressure ventilation | 0 
metabolic derangements | 0 
hemodynamic instability | 0 
vasopressors | 0 
immune response initiation | 0 
complement activation | 0 
thrombin formation | 0 
endothelial inflammation | 0 
non-occlusive mesenteric ischemia | 12 
acute mesenteric ischemia | 12 
small intestinal hypoperfusion | 12 
bowel wall necrosis | 12 
CECT scan showed patent mesenteric vessels | 0 
CECT scan showed collection of fluid | 0 
abdominal X-ray showed multiple air fluid levels | 0 
abdominal X-ray showed prominent dilated small bowel loops | 0 
histopathological report showed small bowel necrosis | 24 
microthrombi in the lamina propria | 24 
microthrombi in the submucosa | 24 
glandular necrosis | 24 
mucosal denudation | 24 
decreased crypts in the lamina propria | 24 
submucosa edematous | 24 
dense acute inflammatory cells | 24 
hyalinized blood vessels | 24 
microthrombi formation | 24 
anticoagulant use | 24 
D-dimer elevated | 0 
fibrinogen elevated | 0 
thromboembolism prophylaxis | 0 
expired | 336 
multi-organ dysfunction syndrome | 168 
Acute Kidney Injury | 168 
sepsis | 168 
reintubation | 144 
COVID pneumonia | 144 
total parenteral nutrition | 24 
low molecular weight Heparin | 24 
Vancomycin IV | 24 
Meropenem IV | 24 
double barrel loop ileostomy | 12 
resection of gangrenous segment | 12 
gangrenous small bowel | 12 
emergency laparotomy | 12 
intravenous antibiotics | 0 
analgesics administered | 0 
supplemental oxygen | 0 
crystalloids administered | 0 
Foley catheterization | 0 
nasogastric tube decompression | 0 
raised lactate level | 0 
metabolic acidosis | 0 
liver function test abnormal | 0 
raised amylase | 0 
leukocytosis | 0 
COVID-19 positive | 0 
sinus rhythm | 0 
tachycardia | 0 
respiratory rate 22 breaths/min | 0 
body temperature 38.7°C | 0 
blood pressure 95/70 mmHg | 0 
oxygen saturation 85% | 0 
vomiting | -72 
palpitation | -72 
abdominal pain aggravated after ingestion of food | -72 
acute abdominal pain | -72 
admitted to the hospital | 0 
female | 0 
57 years old | 0