bilateral otalgia | -120
use of olive oil ear drops | -120
Glasgow Coma Scale score 8 | -120
bilateral green purulent rhinorrhea | 0
bilateral proptosis | 0
right sided chemosis | 0
tachypnoeic | 0
tachycardic | 0
pyrexial | 0
Glasgow Coma Scale score 11 | 0
flexible nasendoscopy | 0
thick green secretions | 0
raised CRP | 1
raised white cell count | 1
raised neutrophil count | 1
low lymphocyte count | 1
raised lactate | 1
pus aspirates collected | 1
Streptococcus pneumoniae isolated | 1
contrast-enhanced computed tomography | 1
opacification of the paranasal sinuses | 1
bony erosion of the lateral walls of both ethmoid sinuses | 1
soft tissue bulging into the right orbit | 1
bilateral proptosis | 1
lumbar puncture | 2
pale cloudy fluid | 2
extremely cellular specimen | 2
high protein | 2
low glucose | 2
Streptococcus pneumoniae isolated | 2
treatment for sepsis and presumed meningitis initiated | 2
intravenous ceftriaxone started | 2
fluticasone nasal spray started | 2
xylometazoline hydrochloride nasal spray started | 2
saline nasal irrigation started | 2
admitted to critical care unit | 3
intubated and ventilated | 12
extubated | 192
completed 10-day course of intravenous antibiotics | 240
discharged home | 312
prescribed betamethasone nasal drops | 312
prescribed fluticasone nasal spray | 312
regular saline nasal irrigation | 312
recovered well | 744
returned to work full time | 744
vivid memories of stay on CCU | 744
no signs of post-traumatic stress disorder | 744
managed medically as an outpatient | 744
contrast-enhanced magnetic resonance imaging | 876
extensive bilateral ethmoid polyposis | 876
hypertrophied inferior turbinates | 876
left sided smooth dural enhancement | 876
Aspergillus and Alternaria specific IgE levels within normal range | 876