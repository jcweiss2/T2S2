18 years old | 0
male | 0
admitted to the emergency department | 0
bite injury to the hand | 0
domesticated animal bite | 0
stray animal bite | 0
human bite | 0
violence-related human bite | 0
clenched fist injury | 0
tooth mark at inoculation site | 0
broken tooth | 0
infection | 0
Eikenella corrodens infection | 0
delayed presentation | 0
Pasteurella infection | 0
tenosynovitis | 0
flexor tenosynovitis | 0
septic arthritis | 0
compartment syndrome | 0
haemorrhagic necrotizing inflammation | 0
paraesthesia | 0
coagulopathy | 0
thrombocytopenia | 0
multiple organ failure | 0
intensive care unit management | 0
blood product substitution | 0
renal support | 0
joint destruction | 0
intra)articular envenomation | 0
popliteal vein thrombosis | 0
complement system activation | 0
amputation of fingers | 0
centipede bite | 0
necrotising fasciitis | 0
cellulitis | 0
severe skin reactions | 0
horse bite | 0
isolated dislocation of the pisiform | 0
marine animal bite | 0
jellyfish sting | 0
median nerve involvement | 0
demyelinating lesion | 0
neuropathic pain | 0
sting ray injury | 0
synovitis | 0
synovectomy | 0
lumbrical muscle necrosis | 0
chronic inflammation | 0
toxic shock syndrome | 0
fish tooth injury | 0
Stonefish envenomation | 0
granulomatous skin lesions | 0
carpal tunnel syndrome | 0
wasp sting | 0
compartment syndrome in child | 0
acute myocardial infarction | 0
lizard bite | 0
ferret bite | 0
Mycobacterium chelonae infection | 0
pyogenic flexor tenosynovitis | 0
osteomyelitis | 0
death due to Capnocytophaga canimorsus septicaemia | 0
external fixation for fractures | 0
patient reported outcome measures | 0
multidisciplinary approach | 0
<|eot_id|>
    