65 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
admitted to the hospital | 0 | 0 | Factual
multiple blisters | -432 | 0 | Factual
erosions | -432 | 0 | Factual
oral mucosa | -432 | 0 | Factual
scalp | -432 | 0 | Factual
superadded maggot infection | -432 | 0 | Factual
previous episodes of lesions | -720 | -168 | Factual
treatment with steroids | -720 | -168 | Factual
unknown generic medications | -720 | -168 | Factual
lesions all over the body | -168 | 0 | Factual
febrile | 0 | 0 | Factual
flaccid blisters | 0 | 0 | Factual
erosions | 0 | 0 | Factual
Nikolsky sign positive | 0 | 0 | Factual
diagnosis of PV | 0 | 0 | Factual
skin biopsy | 0 | 0 | Factual
tzanck smear | 0 | 0 | Factual
intravenous dexamethasone pulse | 0 | 72 | Factual
supportive care | 0 | 72 | Factual
intravenous antibiotics | 0 | 72 | Factual
isolation intensive care unit | 0 | 0 | Factual
oozing from skin ulcerations | 72 | 72 | Factual
hemorrhagic excoriation | 72 | 72 | Factual
peeling of skin | 72 | 72 | Factual
methyl prednisolone | 72 | 168 | Factual
hypoproteinemia | 168 | 168 | Factual
pleural effusion | 168 | 168 | Factual
enterobacter | 168 | 168 | Factual
Staphylococcus aureus | 168 | 168 | Factual
Proteus mirabilis | 168 | 168 | Factual
Tigecycline | 168 | 240 | Factual
vancomycin | 168 | 240 | Factual
sepsis | 168 | 240 | Factual
high grade fever | 168 | 240 | Factual
albumin levels fell | 168 | 240 | Factual
TPE | 240 | 360 | Factual
cyclophosphamide | 360 | 432 | Factual
IV methyl prednisolone | 360 | 432 | Factual
re-epithelization | 360 | 432 | Factual
healing | 432 | 432 | Factual
oral lesions healed | 432 | 432 | Factual
erosions on back | 432 | 432 | Factual
anterior aspect of thigh | 432 | 432 | Factual
buttocks | 432 | 432 | Factual
discharged | 432 | 432 | Factual