80 years old | 0
male | 0
transferred from a peripheral hospital to the university hospital ICU | 0
diagnosed with COVID-19 through bronchoalveolar lavage | 0
intubated | -168
mechanical ventilation | -168
prone positioning | -168
progressive ARDS | 0
multiple organ failure (MOF) | 0
oliguria | 0
septic shock | 0
hepatic dysfunction | 0
mixed acidosis | 0
Sequential Organ Failure Assessment (SOFA) score of 13 | 0
not initiated ECMO | 0
serum creatinine 3.8 mg/dL | 0
potassium 5.9 mmol/L | 0
pH 7.15 | 0
PaCO2 65 mmHg | 0
base excess of -6.6 mmol/L | 0
started on ADVOS device | 0
regional citrate anticoagulation | 0
atrial fibrillation (AF) | 24
digitoxin administered | 24
continuous ultrafiltration performed with ADVOS device | 24
elevated extravascular lung water index (EVLWI) up to 32 mL/kg | 0
normal global end-diastolic volume index (GEDVI) | 0
normal cardiac index (CI) | 0
AF-related increase in GEDVI (827 to 1021 mL/m²) | 24
GEDVI declined from 1021 to 833 mL/m² | 24
elevated PVPI (mean 4.8 ± 1.1) | 0
mean CI 3.1 ± 0.4 mL/min/m² | 0
effective CO2 removal | 0
correction of acidosis | 0
arterial pCO2 69 ± 14 mmHg | 0
post-dialyzer pCO2 27 ± 12 mmHg | 0
CO2 elimination rate 48 ± 23 mL/min | 0
post-dialyzer venous lactate levels lower than pre-dialyzer | 0
acid-base balance controlled | 0
anuria | 0
elevated lactate levels | 0
vasopressor requirement reduced | 24
system clotting | 24
renewed dialysis circuit | 24
improved circulatory parameters after 95 hours of ADVOS | 95
noradrenalin reduced to 0.04 µg/kg/h | 95
Horovitz-Index increased to PaO2/FiO2 116 mmHg | 95
increased driving pressures (22 vs. 18 mbar) | 95
prone-dependent | 95
hemoptysis | 95
positive SARS-CoV-2 PCR | 95
Klebsiella oxytoca detected in tracheal specimens | 95
positive blood cultures | 95
serum and tracheal Aspergillus antigen testing positive | 95
Amphotericin B administered | 95
Meropenem administered | 95
Linezolid administered | 95
increased vasopressor dosage | 95
increased lactate levels | 95
PaO2 85 mmHg | 95
PaO2/FiO2 106 mmHg | 95
PaCO2 38 mmHg | 95
sudden cardiac arrest | 96
coagulopathic and inflammatory parameters increased (D-Dimers 31497 µg/L) | 96
thrombocytopenia (20 109/L) | 96
ferritin up to 15000 µg/L | 96
IL-6 up to 4457 pg/mL | 96
leucocytosis 16 109/L | 96
PCT 4.8 ng/mL | 96
CRP 34 mg/dL | 96
LDH 2967 U/L | 96
GOT 2973 U/L | 96
death | 96
