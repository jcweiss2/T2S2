36 years old | 0
female | 0
admitted to the hospital | 0
pregnancy | 0
IVF performed | -840
previous IVF attempts | -1008
previous mild OHSS | -1008
abdominal enlargement | -720
oocyte retrieval | -720
embryo transfer | -720
human albumin administered | -720
abdominal discomfort | 0
hyperemesis | 0
low urine output | 0
weight gain | 0
distended abdomen | 0
ascites | 0
bilateral pleural effusions | 0
viable intrauterine twin pregnancy | 0
bilateral multiloculated cystic ovaries | 0
increased leukocyte count | 0
thrombocytosis | 0
electrolyte imbalance | 0
elevated liver enzymes | 0
normal thyroid function | 0
elevated serum E2 level | 0
elevated human chorionic gonadotropin level | 0
negative serology for viral hepatitis | 0
OHSS suspected | 0
supportive care initiated | 0
intravenous crystalloid hydration | 0
20% albumin administered | 0
heparin administered | 0
hemoconcentration resolved | 168
discharged to obstetric ward | 168
fever | 168
shivering | 168
renal failure | 168
increased C-reactive protein | 168
respiratory compromise | 168
transvaginal paracentesis | 168
ascitic fluid analysis | 168
Escherichia coli recovered | 168
ceftriaxone initiated | 168
human albumin administered | 168
improved general condition | 216
improved renal function | 216
transvaginal paracentesis repeated | 216
bacteremia documented | 216
Escherichia coli ESBL recovered | 216
piperacillin/tazobactam administered | 216
Acinetobacter baumannii recovered | 216
meropenem administered | 216
discharged from hospital | 1440
readmitted for fetal vitality assessment | 1008
premature rupture of membranes | 1056
Caesarean section performed | 1120
discharged in good condition | 1122