64 years old | 0
    female | 0
    admitted to the hospital | 0
    cough | -360
    fever | -120
    chest tightness | -120
    shortness of breath | -120
    stayed in Wuhan | -408
    returned to Shenzhen | -144
    pharyngeal swab nucleic acid test positive | 0
    COVID-19 diagnosis | 0
    high-flow nasal catheter oxygen therapy | 0
    intermittent noninvasive mechanical ventilation | 0
    interferon atomization | 0
    lopinavir/ritonavir tablets | 0
    gamma globulin | 0
    thymalfasin | 0
    naltrexate calcium | 0
    oxygenation index decreased to 150 mmHg | 120
    invasive mechanical ventilation | 120
    prone position ventilation | 120
    ribavirin | 120
    ceftazidime | 120
    linezolid | 120
    immunoglobulin | 120
    methylprednisolone | 120
    large amount of thin yellow sputum | 168
    CT exudate increased | 168
    CRP increased | 168
    IL-6 increased | 168
    alveolar lavage fluid galactomannan increased | 168
    blood galactomannan increased | 168
    β-glucan level increased | 168
    secondary pulmonary aspergillosis | 168
    voriconazole | 168
    prone position ventilation stopped | 216
    tracheal intubation removed | 240
    nucleic acid test negative | 504
    discharged from ICU | 576
    chest CT resolution of infiltrates | 936
    completely recovered | 936
    discharged | 936
    <|eot_id|>
    