35 years old | 0
male | 0
admitted to the hospital | 0
NYHA Class IV dyspnea | 0
acute pulmonary edema | 0
no hypertension | 0
former smoker | -10080
former morbid obese | -8760
BMI of 26 kg/m2 | 0
previous episode of acute myopericarditis | -5040
fever | -5040
odynophagia | -5040
previous acute pulmonary edema | -5040
admission to the intensive coronary care unit | -5040
echocardiogram showed slightly hypertrophied left ventricle | -5040
ejection fraction of 30% | -5040
akinesia of the interventricular septum | -5040
inferolateral hypokinesia | -5040
no pericardial effusion | -5040
inotropic and depletive treatment | -5040
adequate clinical evolution | -5040
recovered systolic function | -5040
no subsequent cardiac monitoring | -5040
sinus tachycardia | 0
short QRS | 0
repolarization alterations | 0
elevation of the ST segment | 0
ST depression | 0
mild anemia | 0
leukocytosis with left deviation | 0
slight elevation of troponins | 0
acute respiratory acidosis | 0
radiological findings compatible with acute pulmonary edema | 0
moderate left ventricle dysfunction | 0
apical and lateral hypokinesia | 0
intensive depletive treatment | 0
severe hypotension | 2
systolic BP of 60 mmHg | 2
bradycardia | 2
oliguria | 2
vasoactive amines for hemodynamic stabilization | 2
admitted to the Coronary Intensive Care Unit | 2
reversal of systolic dysfunction | 4
reversal of ECG alterations | 4
new echocardiogram | 48
partial recovery of segmental contractility alterations | 48
mild septal hypokinesia | 48
systolic function of 54% | 48
mild left ventricular hypertrophy | 48
moderate dilatation of the left atrium | 48
coronary angiography | 72
no significant coronary abnormalities | 72
cardiac and suprarenal MRI | 72
preserved systolic function | 72
EF 58% | 72
slight inferobasal hypocinesia | 72
solid nodular lesion at the left adrenal gland | 72
pheochromocytoma | 72
delayed enhancement study | 72
subepicardial and inferobasal contrast uptake | 72
myocardial edema | 72
elevated catecholamine excretion | 120
alpha and beta medical blockage | 120
laparoscopic anterior left adrenalectomy | 720
30 mm tumor | 720
no signs of invasion of adjacent structures | 720
postoperative course was favorable | 720
hemodynamically stable | 720
normal tensional controls | 720
discharged | 888
normalized catecholamine excretion | 1008
MRI showed significant decrease of subepicardic enhancement | 1008
preserved ejection function of 63% | 1008
pathology confirmed diagnosis of pheochromocytoma | 1008
no signs of malignancy | 1008