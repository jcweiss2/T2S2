34 years old | 0
male | 0
admitted to intensive care unit | 0
septic shock | 0
multiple organ failure | 0
poor oral intake | 0
fever | 0
altered mental status |9 0
anorexia | 0
dyspnea | 0
alcohol use disorder | 0
no other past medical history | 0
immigrated from Sudan | -70080
employed at meat processing plant | 0
thin | 0
awake | 0
alert | 0
disoriented | 0
scleral icterus | 0
dry mucosal membranes | 0
tachycardia | 0
no murmurs | 0
bilateral rales | 0
rhonchi | 0
soft abdomen | 0
nontender abdomen | 0
distended abdomen | 0
temperature 35.8°C | 0
heart rate 152 bpm | 0
sinus rhythm | 0
respiratory rate 42 breaths per minute | 0
blood pressure 114/75 mmHg | 0
low dose norepinephrine | 0
oxygen saturation 97% | 0
heated high flow nasal cannula oxygen therapy | 0
leukopenia (WBC 2.6 x10³/μL) | 0
elevated lactic acid 4.3 mmol/L | 0
hyperbilirubinemia (total bilirubin 4.3 mg/dL) | 0
direct bilirubin 3.48 mg/dL | 0
elevated AST 423 units/L | 0
elevated ALT 495 units/L | 0
elevated ALP 218 units/L | 0
normal ammonia level | 0
urine toxicology positive for benzodiazepines | 0
acute respiratory acidosis | 0
anion gap metabolic acidosis | 0
hypoxic respiratory failure | 0
COVID-19 PCR positive | 0
microangiopathic hemolytic anemia ruled out | 0
multifocal pneumonia | 0
right-sided pleural effusion | 0
cardiac enlargement | 0
severe hepatosplenomegaly | 0
steatosis | 0
gallstones | 0
pericholecystic fluid | 0
enlarged kidneys | 0
mesenteric edema | 0
diffuse abdominal lymphadenopathy | 0
omental nodularity | 0
dexamethasone treatment for COVID-19 pneumonia | 0
no remdesivir | 0
no tocilizumab | 0
acute hepatic injury | 0
intubation | 24
escalation of antibiotics | 24
worsening renal function | 24
hemodialysis | 24
continued clinical decline | 24
expanded infectious work-up | 24
negative HIV | 24
negative hepatitis B | 24
negative hepatitis C | 24
negative syphilis | 24
negative histoplasma | 24
negative aspergillus | 24
negative cryptococcus | 24
negative candida | 24
negative pneumocystis jirovecii | 24
negative herpes simplex virus 1 | 24
negative herpes simplex virus 2 | 24
negative cytomegalovirus | 24
negative clostridium difficile | 24
negative malaria | 24
Epstein Barr virus past exposure | 24
broad gastrointestinal stool PCR negative | 24
positive sputum cultures (Klebsiella Pneumoniae) | 24
antibiotics de-escalated | 24
positive hepatitis A IgM serology | 24
positive interferon-gamma release assay | 24
latent tuberculosis concern | 24
active tuberculosis diagnosis | 168
dexamethasone discontinued | 24
four-drug TB therapy initiated | 24
TB therapy discontinued | 48
bilirubin increase | 48
rifampin restarted | 72
ethambutol restarted | 72
pyrazinamide restarted | 72
isoniazid held | 24
levofloxacin started | 168
concern for secondary HLH | 168
worsening transaminitis | 168
persistent fever | 168
hepatomegaly | 168
erythropenia | 168
leukopenia | 168
elevated ferritin 77,455.2 ng/ml | 168
elevated triglycerides 252 mg/dl | 168
hypofibrinogenemia 120 mg/dl | 168
elevated CXCL9 232,385 pg/mL | 168
elevated soluble IL-1 receptor alpha 5867 units/mL | 168
bone marrow biopsy deferred | 168
H-score 233 | 168
methylprednisolone initiated | 168
no etoposide | 168
clinical improvement on steroids | 168
tracheostomy | 168
percutaneous endoscopic gastrostomy | 168
recovery of renal function | 168
hemodialysis line removed | 168
discharged to long-term care facility | 216
steroid taper | 216
antituberculosis therapy (rifampin) | 216
antituberculosis therapy (ethambutol) | 216
antituberculosis therapy (pyrazinamide) | 216
antituberculosis therapy (levofloxacin) | 216
