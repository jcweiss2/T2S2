61 years old | 0
male | 0
admitted to the hospital | 0
progressive dyspnoea NYHA class IV | -48
anasarca | -48
ventricular fibrillation | -1464
type 2 amiodarone-induced thyrotoxicosis | -2928
discontinuation of amiodarone | -2928
initiation of thiamazole therapy | -2928
normal thyroid function tests | -48
trans-oesophageal echocardiogram without evidence of intracardiac thrombi | 504
three unsuccessful external defibrillations | 504
re-initiation of oral amiodarone 800 mg/day | 504
discontinuation of amiodarone | 672
acute kidney injury | 1008
anuria | 1008
admission to the intensive care unit | 1008
initiation of continuous veno-venous haemodialysis | 1008
exacerbation of chronic driveline infection | 1032
chronic driveline infection | -7296
post-left ventricular assist device implantation | -52560
clinical deterioration | 1032
shared decision for best supportive care | 1032
death due to septic shock with multi-organ failure | 1104
advanced heart failure | -62640
LVAD support | -62640
dilated cardiomyopathy | -62640
heart failure refractory to medical therapy | -62640
morbid obesity | -62640
body mass index 41 kg/m2 | -62640
arterial pulse absent | 0
normal capillary refill time | 0
normal core temperature | 0
unremarkable neurologic exam | 0
elevated serum creatinine | 0
elevated N-terminal prohormone of brain natriuretic peptide | 0
elevated serum lactate level | 0
global akinesia of all cardiac chambers | 0
profound dilation of the right ventricle | 0
faint movements of the tricuspid valve leaflets | 0
initiation of intravenous furosemide | 0
multiple unsuccessful external defibrillations | 0
initiation of oral amiodarone | 0
severe comorbidities | 0
morbid obesity | 0
severe renal failure | 0
incessant ventricular fibrillation | 0
end-stage renal failure | 24
complications of sepsis | 24
death | 24
