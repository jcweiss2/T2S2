19 years old| 0
    male| 0
    admitted to the emergency department| 0
    fever | -144
    headache | -144
    nausea | -144
    vomiting | -144
    heart rate 134 bpm | 0
    respiratory rate 26 rpm | 0
    blood oxygen saturation 89% | 0
    20,300/mm3 leukocytosis | 0
    16,321/mm3 neutrophils | 0
    58,000/mm3 thrombocytopenia | 0
    431 U/L aspartate transaminase | 0
    145 U/L alanine transaminase | 0
    213.8 mg/L C-reactive protein | 0
    anti-HIV test negative | 0
    renal function unremarkable | 0
    electrolyte levels unremarkable | 0
    brain CT soft tissue enlargement | 0
    extradural collection | 0
    thick content frontal and maxillary sinuses | 0
    sepsis | 0
    admitted to intensive care unit | 0
    sepsis protocol performed | 0
    blood sample collected | 0
    ceftriaxone 2 g every 12 h | 0
    metronidazole 500 mg every 8 h | 0
    oxacillin 2 g every 4 h | 0
    mechanical ventilation needed | 0
    another brain CT scan | 0
    partial sagittal sinus thrombosis | 0
    paranasal sinus CT scan | 0
    right frontal sinus disease | 0
    maxillary sinus disease | 0
    ethmoidal sinus disease | 0
    sinuous nasal septum | 0
    bullous left middle nasal concha | 0
    soft tissue drainage | 24
    neurosurgical drainage | 168
    gram-positive cocci | 0
    anticoagulation initiated | 0
    enoxaparin 40 mg every 12 h | 0
    S. constellatus identified | 0
    resistant to β-lactams | 0
    susceptible to teicoplanin | 0
    susceptible to vancomycin | 0
    anaerobic cultures negative | 0
    no other pathogen identified | 0
    antimicrobial therapy changed | 0
    vancomycin 1.5 g every 12 h | 0
    metronidazole 500 mg every 8 h | 0
    sensory improvement | 672
    no complications | 0
    no adverse reactions | 0
    discharged | 720
    no sequelae at 6-month follow-up | 4320
    
    <|eot_id|>
    