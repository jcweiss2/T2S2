28 years old | 0
female | 0
admitted to the hospital | 0
asymptomatic | 0
large left-to-right shunt | 0
secundum ASD | 0
normal pulmonary venous drainage | 0
normal ventricular function | 0
elevated right atrial pressure | 0
elevated left ventricular end-diastolic pressure | 0
normal pulmonary artery pressure | 0
transcatheter closure | 0
placement of stiff guidewire | 0
delivery sheath in the left upper pulmonary vein | 0
device closure | 0
Cera septal occluder | 0
transesophageal echocardiographic guidance | 0
endotracheal bleeding | 48
protamine | 48
packed red cell transfusion | 48
hemoglobin drop | 48
cardiomegaly | -24
increased pulmonary blood flow | -24
left upper zone infiltrates | 48
lung bleed | 48
progressive respiratory distress | 72
hypoxia | 72
acute respiratory distress syndrome | 72
dilated right heart chambers | 72
biventricular systolic dysfunction | 72
mild pleural effusion | 72
pericardial effusion | 72
elevated right ventricular systolic pressures | 72
pleural effusion | 72
lung collapse | 72
pulmonary edema | 72
elevated inflammatory biomarkers | 72
elevated C-reactive protein | 72
elevated d-Dimer | 72
elevated troponin I | 72
elevated COVID total antibodies | 72
supplemental oxygen | 72
enoxaparin | 72
warfarin | 72
broad-spectrum antibiotic | 72
aspirin | 72
beta-blocker | 72
sildenafil | 72
diuretics | 72
reduction of biomarkers | 120
discharged | 168
hemodynamically stable | 168
asymptomatic | 360
normal effort tolerance | 360
negative RT-PCR for COVID-19 | -24
normal preprocedural blood investigations | -24
COVID-19 infection | -672 
Note: The time stamp is an approximation based on the text and may not be exact. The events that happened before admission have negative timestamps, and the events that happened after admission have positive timestamps. The events with no specific time are assigned a timestamp of 0.