38 years old | 0  
    male | 0  
    admitted to the hospital | 0  
    rectal mucous discharge | -17520  
    family history of pancreatic cancer | 0  
    colonoscopy | -8760  
    nodular-mixed type lateral spreading tumor | -8760  
    histopathology | -8760  
    tubular-villous adenoma with high-grade dysplasia | -8760  
    endorectal ultrasound with 3-dimensional reconstruction | -8760  
    mixed echogenicity image | -8760  
    endoscopic transanal resection | 0  
    no rectal perforation into the peritoneal cavity | 0  
    wound closure with running suture | 0  
    colon mechanical preparation with mannitol | -24  
    surgical antibiotic prophylaxis with ciprofloxacin | -24  
    surgical antibiotic prophylaxis with metronidazole | -24  
    histologic analysis of resected lesion | 0  
    tubular-villous adenoma with high-grade dysplasia | 0  
    intramucosal carcinoma | 0  
    negative surgical margins | 0  
    no abdominal discomfort | 24  
    no nausea | 24  
    no fever | 24  
    tolerance of solid food | 24  
    diffuse abdominal pain | 48  
    asthenia | 48  
    heart rate of 122 beats/min | 48  
    respiratory rate of 25 breaths/min | 48  
    painful abdomen on deep palpation | 48  
    white blood cell count of 10,270/mm3 | 48  
    immature forms 14% | 48  
    serum C-reactive protein level of 25 mg/dL | 48  
    metabolic acidosis | 48  
    elevated lactic acid | 48  
    diagnosis of abdominal focus sepsis | 48  
    volume expansion | 48  
    antibiotics changed to piperacillin-tazobactam | 48  
    admission to intensive care unit | 48  
    abdominal radiography | 48  
    computed tomography of the abdomen with intravenous contrast | 48  
    pneumoretroperitoneum | 48  
    laparotomy | 48  
    diffuse retroperitoneal gas infiltration | 48  
    loop colostomy | 48  
    opening of rectal wound points | 48  
    hospitalization in intensive care unit | 48  
    discharge after 11 days | 264  
    stoma closure after 6 months | 4320  

