28 years old | 0
man | 0
schizophrenia | 0
high-dose clozapine poisoning | 0
admitted to Emergency Department | 0
legal guardian | 0
guardian alerted police | 0
found in apartment | -unknown duration
impaired vigilance | -unknown duration
no physical trauma | -unknown duration
depleted blisters of clozapine (8 g) found | -unknown duration
presumed ingestion of 8 g clozapine | -unknown duration
unclear intent | -unknown duration
no signs of preceding emesis | -unknown duration
somnolent | 0
reduced Glasgow coma scale (11 points) | 0
sinus tachycardia (130/min) | 0
hypertension (157/93 mmHg) | 0
consultation with poisoning center | 0
watch and wait strategy | 0
symptomatic therapy | 0
cranial CT | 0
no cerebral pathologies | 0
thoracic CT | 0
pulmonary infiltrates | 0
atelectasis | 0
pneumomediastinum | 0
soft-tissue emphysema | 0
rhabdomyolysis | 0
crush syndrome | 0
acute renal failure AKIN II | 0
creatinine (188 µmol/l) | 0
myoglobin (6231 µg/l) | 0
creatine kinase (367 µkat/l) | 0
urine investigations | 0
no evidence of other drugs | 0
progressive impairment of vigilance | 0
respiratory insufficiency | 0
GCS=7 | 0
peripheral oxygen saturation < 90% | 0
respiratory rate 26/min | 0
invasive ventilation | 0
no fever | 0
bronchoscopy | 0
esophagogastroduodenoscopy | 0
no anatomical air leakage | 0
SOFA score 15 | 0
sepsis | 0
community-acquired bilateral pneumonia | 0
treated with Piperacillin/Tazobactam | 0
admitted to ICU | 10
septic shock | 10
required vasopressors | 10
vasopressors tapered after fluid supplementation | 10
hypertension | 10
moderate tachycardia | 10
sodium nitroprusside required | 10
successful respiratory weaning | 31
extubated | 31
respiration remained stable | 31
drowsiness (Richmond Agitation-Sedation Scale -2) | 31
tachycardia | 31
hypertension | 31
inadequate communication | 31
hyposalivation | 31
anticholinergic syndrome | 31
treated with physostigmine | 31
became more awake (Richmond Agitation-Sedation Scale 0) | 31
tachycardia resolved | 31
hypertension resolved | 31
physostigmine therapy stopped | after 2 days (48 hours)
follow-up CT at day 6 | 144
pneumomediastinum regressed | 144
soft-tissue emphysema regressed | 144
pneumonia in healing process | 144
serum clozapine levels decreased to therapeutic at day 4 | 96
transferred to Psychiatry Department | 144
confirmed clozapine intake | 144
denied suicidal intention | 144
completely awake (Richmond Agitation-Sedation Scale 0) | 144
oriented | 144
good general condition | 144
good respiratory condition | 144
no oxygen needed | 144
regression of renal failure | 144
regression of rhabdomyolysis | 144
regression of inflammation | 144
creatinine (78 µmol/l) | 144
myoglobin (145 µg/l) | 144
white blood count (10.5 GPt/l) | 144
