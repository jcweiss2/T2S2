26 years old | 0
male | 0
admitted to the hospital | 0
restrictive subaortic VSD | -2160
mild pulmonary hypertension | -2160
hypochromic anemia | -2160
fatigue | -2160
effort limitation | -2160
exertional dyspnea | -2160
ascites | -2160
persistent inflammatory syndrome | -2160
weight loss | -2160
increased blood cell count | 0
C-reactive protein | 0
procalcitonin | 0
anemia | 0
thrombocytopenia | 0
echocardiography | 0
IE with mobile vegetations | 0
severe regurgitation of the aortic valve | 0
severe regurgitation of the tricuspid valve | 0
severe regurgitation of the pulmonary valve | 0
aortic annulus abscess | 0
severe biventricular dysfunction | 0
severe PHT | 0
septic shock | 0
multiple organ dysfunction syndrome | 0
hypotensive | 0
hypoxemic | 0
severe metabolic acidosis | 0
oliguria | 0
neurologic dysfunction | 0
mechanical ventilation | 0
hemodynamic support | 0
dobutamine | 0
norepinephrine | 0
continuous venovenous hemodiafiltration | 0
cytokine removal filter | 0
Gram-negative bacilli | 0
meropenem | 0
clinical improvement | 168
weaning of norepinephrine | 168
weaning of mechanical ventilation | 168
organ functions recovered | 168
ventricular function improved | 168
paroxysmal supraventricular tachycardia | 384
septic discharge | 384
recurrence of septic shock | 384
hemodynamic deterioration | 384
lactate increase | 384
transient hepatic cytolysis | 384
oliguria | 384
electrical conversion | 384
administration of dobutamine | 384
administration of levosimendan | 384
surgery | 432
bicaval-aortic cardiopulmonary bypass | 432
Custodiol cardioplegia | 432
aortic valve replacement | 432
tricuspid valve replacement | 432
pulmonary valve replacement | 432
aortic annulus abscess debridement | 432
VSD closure | 432
postoperative outcome | 456
stable hemodynamics | 456
no arrhythmias | 456
extubation | 456
Milrinone infusion | 456
inotrope withdrawal | 480
sacubitril/valsartan treatment | 480
discharge | 720
follow-up | 4320
resumed work | 4320
normally functioning valves | 4320
improved ventricular function | 4320
no sign of infection | 4320
follow-up | 7776
asymptomatic | 7776
sacubitril/valsartan treatment | 7776
LVEF | 7776