39 years old | 0
female | 0
palpable mass on her right breast | -168
Hodgkin lymphoma | -6336
chemotherapy | -6336
mantle field radiation | -6336
inflammatory colitis | -6336
mesalazine | -336
family history of myxoid liposarcoma | 0
breast radiological examination | -168
invasive ductal carcinoma | -168
triple-negative phenotype | -168
MIB1 85% | -168
staging CT scan | -168
neoadjuvant chemotherapy | -112
paclitaxel | -112
carboplatin | -112
port-à-cath insertion | -84
subcutaneous cellulitis | -60
colliquative necrosis | -60
fever | -60
elevated white blood cell count | -60
neutrophilia | -60
elevated C-reactive protein | -60
broad-spectrum i.v. antibiotic therapy | -60
piperacillin/tazobactam | -60
daptomycin | -60
PORT rimotion | -60
necrosectomy | -60
defervescence | -54
improvement in subcutaneous cellulitis | -54
febrile seizure | -48
WBC rise | -48
worsening of skin lesion | -48
second necrosectomy | -48
peripheral blood cultures | -48
skin plug | -48
i.v. catheter tip positivity for Klebsiella pneumoniae | -48
antibiotic therapy modification | -48
meropenem | -48
levofloxacin | -48
chest/abdomen CT scan | -48
mediastinitis | -48
bilateral pleural effusion | -48
left pulmonary atelectasis | -48
thoracoscopy | -42
pleural and mediastinal drainage | -42
sepsis | -42
broad-spectrum antibiotic and antifungal therapy | -42
hemodynamic support | -42
non-invasive ventilation | -42
specimens of skin and subcutaneous and muscular tissue analysis | -42
intensive inflammatory infiltrate | -42
neutrophils | -42
systemic methylprednisolone | -24
topical cyclosporine | -24
seriate chest X-ray | -24
CT scan | -24
progressive resolution of mediastinitis | -24
progressive resolution of pleural effusion | -24
wound improvement | -24
scar | -24
blood works normalization | -24
breast ultrasound | -12
no change in the dimension of the lump | -12
multidisciplinary meeting | -12
right mastectomy | 0
axillary dissection | 0
breast surgical wound healing | 12
pathology assessment | 12
fibroelastosis | 12
chronic inflammation | 12
isolated neoplastic cells | 12
negative axillary nodes | 12
restaging brain/chest/abdomen CT | 12
negative for distant metastasis | 12
BRCA and p53 mutation tests | 12
negative | 12
autologous skin graft | 24
no further complications | 24
PICC implant | 24
chemotherapy with carboplatin and paclitaxel | 24
dose reduction | 24
good tolerance | 168
follow-up | 168