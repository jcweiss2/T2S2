64 years old | 0
female | 0
Hepatitis C-induced liver cirrhosis | -8760
end-stage renal disease | -8760
hemodialysis | -8760
chronic anemia | -8760
hypothyroidism | -8760
admitted to the emergency department | 0
fatigue | -72
weakness | -72
blurry vision | -72
shortness of breath | -72
fishing in a pond | -72
fell | -72
abrasion on her left forearm | -72
blisters on her left forearm | -24
blood pressure 60/26 mmHg | 0
pulse rate 88/min | 0
respiration rate 17/min | 0
T 94.0 F | 0
hyperpigmentation | 0
edema | 0
hemorrhagic bullae | 0
diminished breath sounds | 0
bibasilar crackles | 0
white blood cell count 19,550 | 0
lactic acid 10.7 mmol/L | 0
bibasilar atelectasis | 0
consolidation consistent with pneumonia | 0
hepatosplenomegaly | 0
portal venous hypertension | 0
ascites | 0
septic shock | 0
cellulitis | 0
pneumonia | 0
pressors | 0
admitted to the intensive care unit | 0
Infectious disease consultations | 0
Aeromonas infection suspected | 0
gentamicin | 0
Levaquin | 0
vancomycin | 0
Zosyn | 0
orthopedic surgery consulted | 0
blisters aspirated | 24
no excisional debridement | 24
white blood cell count 12,350 | 48
blood cultures released | 72
Aeromonas veronii complex | 72
ampicillin-sulbactam resistant | 72
piperacillin-tazobactam resistant | 72
antibiotics narrowed down | 96
post-dialysis ceftazidime | 96
gentamicin | 96
post-dialysis vancomycin | 96
discharged | 240