79 years old | 0
    woman | 0
    admitted to the emergency department | 0
    fever | -120
    malaise | -120
    anorexia | -120
    confusion | -96
    unconsciousness | -96
    diabetes (type 2 diabetes) | 0
    hypertension | 0
    atrial fibrillation | 0
    cholecystectomy | 0
    appendectomy | 0
    pyrexia (maximum temperature 39°C) | 0
    noninvasive mechanical ventilation | 0
    normal blood pressure (120/90 mmHg) | 0
    tachycardia (155 bpm) | 0
    indifferent attitude | 0
    decreased breath sounds | 0
    soft abdomen | 0
    no peripheral edema | 0
    increased procalcitonin level (31 ng/mL) | 0
    high white blood cell count (12.21 × 10⁹/L) | 0
    anemia (hemoglobin 93 g/L) | 0
    low platelet cell count (22 × 10⁹/L) | 0
    elevated NT-pro-BNP levels (14100 pg/mL) | 0
    abdominal US showed non-homogeneous echo zone in left liver lobe | 0
    gas bubbles in hepatic vein | 0
    gas bubbles in inferior vena cava | 0
    gas bubbles in right atrium | 0
    no abnormal hepatic artery perfusion | 0
    no abnormalities in echocardiography | 0
    poor CT image quality due to inability to hold breath | 0
    CT showed irregularly mixed lower-density lesions in liver | 0
    gas density inside liver lesions | 0
    small gas density in adjacent liver parenchyma | 0
    CT report indicated ruptured liver abscess | 0
    CT report indicated intrahepatic bile duct pneumatosis | 0
    blood cultures grew K. pneumoniae | 0
    diagnosed with ruptured K. pneumoniae liver abscess leading to HVG | 0
    administered imipenem and cilastatin | 0
    infection index improvement | 0
    treatment changed to cefoperazone sulbactam | 0
    general supportive measures | 0
    no specific treatment for HVG formation | 0
    gradual improvement | 0
    bedside US revealed no further gas in hepatic vein | 48
    bedside US revealed no further gas in liver abscess | 48
    small liquefaction zone in abscess area | 48
    subsequent follow-up US examinations | 0
    abscess shrank and disappeared | 0
    no other abscess formation | 0
    discharged after 41 days of treatment | 984
    