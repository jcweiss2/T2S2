20 years old | 0
female | 0
admitted to the emergency room | 0
signs of sepsis | 0
hypotension | 0
multi-organ failure | 0
insulin-dependent diabetes mellitus | -672
pulmonary tuberculosis | -144
productive cough | -720
weight loss | -720
fever | -720
anti-tuberculous medicines | -144
CT scan | 0
multiple cavitatory lesions in the right lung | 0
moved to the intensive care unit | 0
insulin infusion | 0
diabetic ketoacidosis | 0
hypoxia | 2
acidosis | 2
pulseless ventricular tachycardia | 2
advance cardiac life support | 2
intubated | 2
endotracheal tube | 2
operating room | 4
VATS | 4
evacuation of the abscess | 4
clinical monitoring | 4
ECG | 4
End-tidal CO2 | 4
pulse oximeter | 4
central venous pressure | 4
invasive blood pressure | 4
anesthesia machine | 4
Isoflurane | 4
FiO2 | 4
air | 4
oxygen | 4
nitrous oxide | 4
left lateral | 4
cis-atracurium | 4
morphine | 4
evacuation of the abscess | 4
major air leak | 6
hypoxia | 6
jet ventilation | 6
Sander's Manu jet Ventilator | 6
ruptured lung abscess | 6
right upper lobe | 6
lung isolation | 8
left sided 32Fr Mallinckrodt double lumen tube | 8
C-Mac Video Laryngoscope | 8
tracheal lumen | 8
clamped | 8
left lung | 8
ventilated differentially | 8
recruitment maneuver | 10
oxygen saturation | 10
right upper lobe lobectomy | 12
packed red blood cell | 12
transfused | 12
phenylephrine | 12
hypotension | 12
boluses | 12
wound closed | 14
chest drain | 14
double-lumen endotracheal tube | 14
single lumen PVC tube | 14
video laryngoscope | 14
ICU | 14
stable condition | 14
bronchoscopy | 24
stump site | 24
no residual defect | 24
discharged | 48