65 years old | 0
female | 0
obesity | 0
type 2 diabetes mellitus | 0
hypertension | 0
hyperlipidaemia | 0
transient ischaemic attack | 0
left-sided breast cancer | 0
fever | -168
dry cough | -168
exertional dyspnoea | -168
hypoxia | -3
bilateral lung ground-glass opacities | -3
SARS-CoV-2 positivity | -3
admitted to the hospital | 0
aspirin | 0
losartan-hydrochlorothiazide | 0
simvastatin | 0
levothyroxine | 0
omeprazole | 0
metformin | 0
liraglutide | 0
diminished breath sounds | 0
bilateral infiltrates | 0
pneumonitis | 0
remdesivir | 0
ceftriaxone | 0
azithromycin | 0
community-acquired pneumonia | 0
acute biventricular heart failure | 168
acute respiratory distress syndrome | 168
acute kidney injury | 168
ischaemic hepatitis | 168
cytokine storm | 168
rapid-sequence intubation | 168
transfer to the medical intensive care unit | 168
tocilizumab | 176
norepinephrine | 176
vasopressin | 176
dobutamine | 176
sodium bicarbonate | 176
inhaled epoprostenol | 176
hydrocortisone | 176
propofol | 176
fentanyl | 176
cisatracurium | 176
clinical improvement | 200
down-trending inflammatory markers | 200
titration off norepinephrine | 200
titration off vasopressin | 200
titration off dobutamine | 200
titration off sodium bicarbonate | 200
cessation of neuromuscular blockade | 200
myocardial recovery | 216
LVEF of 64% | 216
mild RV dysfunction | 216
Grade 2 diastolic dysfunction | 216
small circumferential pericardial effusion | 216
tracheostomy | 240
discharge from the ICU | 240
discharge from the hospital | 336