79 years old | 0
man | 0
German descent | 0
sudden-onset abdominal pain | 0
collapsed | 0
pale | 0
hypotensive | 0
blood pressure 65/40 mmHg | 0
bradycardic | 0
heart rate 40 to 50 beats/minute | 0
slow atrial fibrillation | 0
open exploratory laparotomy | 0
ruptured infrarenal abdominal aortic aneurysm | 0
open repair of aneurysm | 0
significant blood loss | 0
cell saver returning 5.5 L of blood | 0
received 6 units of packed cells | 0
received 4 units of fresh-frozen plasma | 0
received 6 units of cryoprecipitate | 0
received 1 pooled bag of platelets | 0
received 4 L of crystalloids | 0
postoperative intensive care unit admission | 0
intubated | 0
requiring high dose of vasopressors | 0
repeated transthoracic echocardiography | 0
normally functioning heart | 0
no significant ventricular or valvular abnormality | 0
hypertension | -infinity (preexisting condition, timestamp assigned as negative infinity as prior to admission)
benign prostatic hypertrophy | -infinity (preexisting condition, timestamp assigned as negative infinity as prior to admission)
atorvastatin | -infinity (prior to admission)
amlodipine | -infinity (prior to admission)
dutasteride-tamsulosin | -infinity (prior to admission)
allergy to penicillin | -infinity (prior to admission)
rash | -infinity (prior to admission)
postoperative instability | 0
acute kidney injury | 0
mild abdominal hypertension | 0
requiring sedation | 0
requiring paralysis | 0
did not tolerate enteral feeding | 0
received full total parenteral nutrition | 0
extubated | 240 (postoperative day 10)
re-intubated | 240 (a few hours later)
worsening respiratory failure | 240
signs of sepsis | 240
fever | 240
leukocytosis | 240
later became unstable | 240
required vasopressors | 240
source of infection unclear | 240
meropenem commenced | 240
vancomycin commenced | 240
Serratia marcescens isolated in blood cultures | 240
sensitive to meropenem, ciprofloxacin, co-trimoxazole | 240
resistant to penicillins and cephalosporins | 240
Serratia marcescens isolated in urine cultures | 240
Serratia marcescens isolated in sputum cultures | 240
Serratia marcescens isolated in wound swab culture | 264 (2 days later)
hemodynamic improvement | 264
renal function improvement | 264
ventilator-dependent | 264
encephalopathic | 264
tracheostomy | 336 (postoperative day 14)
hyperbilirubinemia | 336
mildly deranged liver transaminase levels | 336
biochemical markers of cholestasis | 336
attributed to bile duct obstruction | 336
no evidence of cholelithiasis | 336
no dilation of biliary ducts | 336
bilirubin continued to increase to 200 µmol/L | 336
ERCP performed | 336
transcutaneous hepatic cholangiography performed | 336
patent right and left hepatic ducts | 336
patent common biliary ducts | 336
smooth tapering toward ampulla | 336
patent cystic duct | 336
stent inserted in common bile duct | 336
8.5-French external biliary drain inserted | 336
no improvement following cholangiography | 336
external biliary drain producing 600 mL of bile | 336
direct bilirubin 300 µmol/L | 432 (postoperative day 18)
conjugated bilirubin 169 µmol/L | 432
repeated abdominal CT showed no intra-abdominal collection | 432
no evidence of bleeding | 432
no other new pathology | 432
subsequent cholangiogram | 432
stent and bile ducts remain patent | 432
meropenem changed to ciprofloxacin | 432
suspicion of VBDS | 432
decrease in bilirubin level | 432
meropenem restarted | 504 (postoperative day 21)
worsening fever | 504
worsening sepsis | 504
increase in serum bilirubin level | 504
meropenem-induced VBDS suspected | 504
antibiotic therapy changed to ciprofloxacin and metronidazole | 552 (postoperative day 23)
dramatic decrease in bilirubin level | 552
bilirubin normalized | 552
clindamycin | 24 (POD1-3)
meropenem | 240 (POD10-18), 504 (POD21-23)
metronidazole | 552 (POD23-38)
ciprofloxacin | 552 (from POD23 to discharge)
vancomycin | 240 (POD10-15)
paracetamol | 24 (POD1-5)
other medications (sedation, analgesia, TPN) | 0 (continuous during admission)
biliary drain plugged | 720 (after 3 days from postoperative day 18)
biliary drain removed | 720
prolonged ICU stay | 720
ventilator-dependent | 720
gradually improved | 720
decannulated | 720
discharged from ICU | 2160 (3-month stay)
no significant organ dysfunction | 2160
treated in general ward | 2160
discharged from hospital | 2160 (final discharge)
