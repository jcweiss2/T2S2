17 years old | 0
female | 0
admitted to the hospital | 0
acute onset of behavioral change | 0
extreme politeness | 0
obedience | 0
pre-morbid gregarious personality | -672
progression to excessive and irrelevant talks | -672
features of disinhibition | -672
frank psychotic features | -240
verbal aggression | -240
physical aggression | -240
muttering to herself | -240
marked delusional thoughts | -240
tendency to run amok | -240
diagnosis of acute functional psychosis | -240
oleanzapine started | -240
behavioral syndrome persisted | -240
mild reduction of psychomotor activity | -240
stiffness of whole body | -240
akinesia | -240
mutism | -240
evaluated by neurologist and psychiatrist | -240
MRI brain scattered T2 and FLAIR hyperintensities | -240
CSF examination no cells | -240
normal CSF protein | -240
normal CSF glucose levels | -240
negative CSF viral markers | -240
negative VDRL test | -240
negative gram stain | -240
negative AFB stain | -240
negative India ink | -240
negative cryptococcal antigen | -240
negative bacterial cultures | -240
negative mycobacterial cultures | -240
negative fungal cultures | -240
EEG non-specific diffuse theta delta slowing | -240
low grade fever | -240
serum Creatinine Phosphokinase raised to 1800 U/dl | -240
diagnosis of NMS due to oleanzapine | -240
dantrolene started | -240
hydration started | -240
slight reduction of rigidity | -240
no other improvement noticed | -240
clinical worsening over next 2 weeks | 336
increasing mental obtundation | 336
persistent akinetic mute state | 336
frequent bouts of tachypnea | 672
tachycardia | 672
hypotension | 672
sweating | 672
deterioration over next 48 hours | 720
gasping for breath | 720
oxygen desaturation | 720
endotracheal intubation | 720
mechanical ventilation | 720
brought to our center | 720
widely fluctuating heart rate | 720
widely fluctuating blood pressure | 720
stimulus-induced sinus tachycardia | 720
tachypnea | 720
diaphoresis | 720
sedative infusion | 720
provisional diagnosis of sepsis syndrome | 720
bilateral aspiration pneumonia | 720
received critical care | 720
received medical support | 720
re-evaluated by neurology team | 720
possibility of immune encephalitis considered | 720
MRI brain repeated | 720
similar changes as before | 720
normal infectious meningoencephalitis workup | 720
CSF samples sent for anti-NMDA receptor antibody | 720
CSF samples sent for anti-VGKC antibody | 720
