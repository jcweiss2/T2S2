56 years old | 0
    man | 0
    presented to the emergency department | 0
    increasing dyspnea | -336
    productive cough | -336
    blood pressure 127/93 mm Hg | 0
    heart rate 99 beats/min | 0
    temperature 86.6°F | 0
    respiratory rate 28/min | 0
    97% saturation on 2L O2 by nasal cannula | 0
    anxious | 0
    jugular venous distention | 0
    bilateral rales | 0
    wheezing | 0
    regular cardiac rhythm | 0
    no evident murmurs | 0
    no S3 | 0
    no S4 | 0
    left lower extremity below the knee amputation | 0
    right lower extremity with 1+ pitting edema | 0
    acute decompensated congestive heart failure | 0
    decompensated chronic pulmonary disease | 0
    furosemide 80 mg IV | 0
    nebulized bronchodilator therapy | 0
    methylprednisolone 125 mg IV | 0
    respiratory status rapidly declined | 0
    admitted to the intensive care unit | 0
    bilevel positive airway pressure | 0
    additional treatment | 0
    developed shock | 0
    multisystem organ failure | 0
    hypoxemic respiratory failure | 0
    hypercapnic respiratory failure | 0
    refractory to BiPAP | 0
    intubated | 0
    vasopressor therapy | 0
    nonischemic cardiomyopathy | 0
    left ventricular ejection fraction of 20%-25% | 0
    status post biventricular implantable cardioverter defibrillator | 0
    status post 25 mm CarboMedics bi-leaflet mechanical aortic valve | 0
    paroxysmal atrial fibrillation | 0
    warfarin | 0
    intermittent noncompliance | 0
    labile INR values | 0
    chronic hypertension | 0
    hyperlipidemia | 0
    tobacco abuse | 0
    ongoing 1.5 ppd use | 0
    chronic kidney disease stage IIIb | 0
    non-insulin-dependent diabetes mellitus | 0
    major depressive disorder | 0
    history of psychotic features | 0
    suicidal ideation | 0
    recurrent noncompliance with medical therapy | 0
    acute decompensated heart failure | 0
    pulmonary thromboembolism | 0
    decompensated chronic pulmonary disease with cor pulmonale | 0
    septic shock | 0
    prosthetic valve dysfunction | 0
    infectious endocarditis | 0
    acute coronary syndrome | 0
    transthoracic echocardiogram | 0
    mechanical aortic valve stenosis | 0
    peak velocity of 4.7 m/s | 0
    acceleration time of 110 ms | 0
    mean gradient of 52 mm Hg | 0
    Doppler velocity index of 0.25 | 0
    mild aortic regurgitation | 0
    Swan-Ganz placement | 0
    intra-aortic balloon pump insertion | 0
    fluoroscopy of the mechanical aortic valve | 0
    fixed nonmobile leaflet | 0
    presumed thrombosis | 0
    history of medication noncompliance | 0
    prohibitively high surgical risk | 0
    alteplase 10 mg IV bolus | 0
    alteplase 90 mg IV infusion over 20 h | 0
    adjuvant therapeutic anticoagulation with heparin infusion | 0
    aPTT at 1.5-2.0 times control value | 0
    serial transthoracic echocardiograms over 4 days | 96
    improvement of mechanical aortic valve function | 96
    peak velocity of 3.6 m/s | 96
    mean pressure gradient of 35 mm Hg | 96
    repeat fluoroscopic evaluation | 96
    normal bi-leaflet motion | 96
    successful thrombolysis | 96
    restoration of function | 96
    no major bleeding events | 96
    no complications | 96
    continued to improve | 96
    successfully extubated | 96
    discharged | 96
    strict instructions to comply with warfarin therapy | 96
    follow-up transthoracic echocardiogram 3 months later | 2160
    normal functioning mechanical aortic valve | 2160
    peak velocity of 2.3 m/s | 2160
    mean pressure gradient of 11 mm Hg | 2160
    <|eot_id|>