49 years old | 0
female | 0
wheelchair-bound | 0
multiple sclerosis | 0
natalizumab treatment | -672
presented to the intensive care unit | 0
prolonged encephalopathy | 0
breakthrough seizures | 0
hypothermia | 0
hypotension | 0
tachycardia | 0
tachypnea | 0
hypoxia requiring mechanical ventilation | 0
elevated white blood cell count | 0
hemoglobin 10.0 g/dL | 0
platelet count 511,000/uL | 0
urine toxicology screen unrevealing | 0
encephalopathy thought to be toxic metabolic cause secondary to sepsis due to pneumonia | 0
started on cefepime | 0
started on vancomycin | 0
continuous EEG monitoring | 0
no seizure activity | 0
antiepileptic medication dosing adjusted | 0
mental status unchanged | 0
MRI brain with contrast | 0
lumbar puncture | 0
MRI showed symmetric marked edema bilateral basal ganglia | 0
mass effect on lateral ventricles | 0
CSF lymphocytic pleocytosis 95 cells/uL | 0
low CSF glucose 29 mg/dL | 0
high protein 103.1 mg/dL | 0
consistent with viral encephalitis | 0
JC virus testing negative | 0
other viral studies negative | 0
viral PCR positive for herpes encephalitis type 2 | 0
started on intravenous acyclovir | 0
improvement in mental status | 0
discharged to rehabilitation center | 0
fever | -72
headache | -72
altered mental status | -72
nausea | -72
vomiting | -72
receptive aphasia | -72
hemiparesis | -72
seizures | -72
meningeal signs | -72
pneumonia | -72
sepsis | -72
natalizumab discontinued | -672
herpes encephalitis type 2 | 0
