61 years old | 0
    male | 0
    admitted to the hospital | 0
    intermittent high-grade fever | -720
    swelling of right knee joint | -720
    severe pain (right knee) | -720
    inability to weight bear | -720
    inability to walk due to knee pain | -168
    urinary tract infection | -720
    type II diabetes mellitus | -720
    sudden onset breathlessness | -24
    emergency department arrival | 0
    consciousness | 0
    febrile | 0
    tachycardic | 0
    tachypnoeic | 0
    hypotensive | 0
    reduced saturation | 0
    extensive bilateral crepitations | 0
    right knee swelling (warm and tender) | 0
    septic arthritis right knee | 0
    severe septicemia | 0
    septic shock | 0
    intubation | 0
    fluid resuscitation | 0
    inotropes administration | 0
    vasopressors administration | 0
    transfer to critical care unit | 0
    intravenous meropenem | 0
    intravenous teicoplanin | 0
    blood gas analysis revealing severe metabolic acidosis | 0
    lactic acidemia | 0
    anuria | 0
    severe leukopenia | 0
    deranged liver function | 0
    deranged renal function | 0
    deranged coagulation profile | 0
    ventricular tachycardia | 0
    cardioverted | 0
    bradycardia | 0
    cardiopulmonary resuscitation (3 cycles) | 0
    death | 24
    blood culture taken | 0
    Gram-negative organism identification | 12
    Burkholderia pseudomallei confirmation | 12
    resistant to polymyxin B | 12
    resistant to aminoglycosides | 12
    susceptible to ceftazidime | 12
    susceptible to co-trimoxazole | 12
    susceptible to carbapenems | 12
    meropenem administration | 0
    teicoplanin administration | 0
    septic shock | 0
    hemodynamic instability | 0
    broad-spectrum antibiotics history | -720

    <|eot_id|>
    61 years old | 0
male | 0
admitted to the hospital | 0
intermittent high-grade fever | -720
swelling of right knee joint | -720
severe pain (right knee) | -720
inability to weight bear | -720
inability to walk due to knee pain | -168
urinary tract infection | -720
type II diabetes mellitus | -720
sudden onset breathlessness | -24
emergency department arrival | 0
consciousness | 0
febrile | 0
tachycardic | 0
tachypnoeic | 0
hypotensive | 0
reduced saturation | 0
extensive bilateral crepitations |5
right knee swelling (warm and tender) | 0
septic arthritis right knee | 0
severe septicemia | 0
septic shock | 0
intubation | 0
fluid resuscitation | 0
inotropes administration | 0
vasopressors administration | 0
transfer to critical care unit | 0
intravenous meropenem | 0
intravenous teicoplanin | 0
blood gas analysis revealing severe metabolic acidosis | 0
lactic acidemia | 0
anuria | 0
severe leukopenia | 0
deranged liver function | 0
deranged renal function | 0
deranged coagulation profile | 0
ventricular tachycardia | 0
cardioverted | 0
bradycardia | 0
cardiopulmonary resuscitation (3 cycles) | 0
death | 24
blood culture taken | 0
Gram-negative organism identification | 12
Burkholderia pseudomallei confirmation | 12
resistant to polymyxin B | 12
resistant to aminoglycosides | 12
susceptible to ceftazidime | 12
susceptible to co-trimoxazole | 12
susceptible to carbapenems | 12
meropenem administration | 0
teicoplanin administration | 0
septic shock | 0
hemodynamic instability | 0
broad-spectrum antibiotics history | -720