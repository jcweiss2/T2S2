40 years old | 0
African-American | 0
female | 0
history of chronic eczema | -672
history of alcohol abuse | -672
history of gout | -672
history of hypothyroidism | -672
worsening eruption | 0
intermittent diarrhea | 0
desquamation of the hands | -336
desquamation of the feet | -336
desquamation of the perioral skin | -336
desquamation of the perineal skin | -336
pain | -336
swelling | -336
hair loss | -336
increasing weakness | -336
fatigue | -336
unintentional weight loss | -336
70 pounds of unintentional weight loss | -336
1 to 2 glasses of wine a day | -336
smoking | -336
erythematous desquamative patches | 0
erosions | 0
crusted lesions | 0
diffuse nonscarring alopecia | 0
scaling patches on the vermillion lips | 0
methicillin-resistant Staphylococcus aureus sepsis | 0
Escherichia coli sepsis | 0
pneumonia | 0
ventilator respiratory support | 0
systemic antibiotics | 0
low zinc levels | 0
positive antitransglutaminase antibodies | 0
positive antiendomysium antibodies | 0
focal villi blunting | 0
Brunner's gland hyperplasia | 0
gluten-free diet | 0
zinc sulfate | 0
resolution of gastrointestinal symptoms | 96
resolution of cutaneous symptoms | 96