28 weeks of gestational age | 0  
    male | 0  
    premature | 0  
    very-low-birth-weight | 0  
    bloody stools | 0  
    NEC (stage 3A) | 0  
    increased gastric residual | -24  
    apnoea | -24  
    grossly bloody stools | -24  
    abdominal distention | -24  
    left abdominal tenderness | -24  
    sluggish bowel sounds | -24  
    increased CRP levels | -24  
    decreased WBC levels | -24  
    positive stool occult blood | -24  
    pneumatosis intestinalis | -24  
    pale | -24  
    less active | -24  
    tachycardia | -24  
    hypotension | -24  
    conventional mechanical ventilation | -24  
    fluid resuscitation | -24  
    haemodynamic support | -24  
    IV antibiotics (piperacillin/tazobactam and vancomycin) | -24  
    E. coli positive blood culture | -96  
    IV antibiotics changed to piperacillin/tazobactam and meropenem | -96  
    clinical improvement | -168  
    radiological improvement | -168  
    resumed EBM feedings | -168  
    second episode of bloody stools | -696  
    soft abdomen | -696  
    non-tender abdomen | -696  
    active bowel sounds | -696  
    positive stool occult blood | -696  
    normal CRP levels | -696  
    normal WBC levels | -696  
    mild thickening of the small bowel | -696  
    no pneumatosis intestinalis | -696  
    antibiotic therapy | -696  
    suspended feeding | -696  
    normal CRP levels | -744  
    normal WBC levels | -744  
    resumed enteral feeding with breast milk | -744  
    negative blood culture | -744  
    third episode of bloody stools | -1104  
    no emesis | -1104  
    no abdominal distension | -1104  
    active bowel sounds | -1104  
    decreased WBC levels | -1104  
    normal CRP levels | -1104  
    mild increase in eosinophil counts | -1104  
    suspected FPIES | -1104  
    suspended feeding | -1104  
    symptoms disappeared | -1104  
    resumed expressed mother's milk without cow's milk | -1104  
    fourth episode of bloody stools | -1296  
    abdominal distension | -1296  
    grossly bloody stools | -1296  
    normal WBC levels | -1296  
    normal CRP levels | -1296  
    increased eosinophil count (13.8%) | -1296  
    suspected FPIES | -1296  
    changed to hydrolyzed formula | -1296  
    resolution of symptoms | -1296  
    diagnosed with FPIES | 0  
    discharged home | 1440  
    nonrecurrence of symptoms | 1440  
    breastfed for 8 months | 1440  
    no bloody stools recurrence | 1440  

