76 years old | 0
    woman | 0
    presented to the Department of Endocrinology, Peking University International Hospital | 0
    progressive neck pain | -720
    neck pain exacerbated by swallowing | -720
    productive cough with yellow sputum | -720
    denied fever | 0
    denied weight loss | 0
    II° thyroid enlargement | 0
    indurated texture | 0
    no thyroid bruits | 0
    lungs clear to auscultation bilaterally | 0
    no dry rales | 0
    no wet rales | 0
    pre-hospital thyroid function tests | 0
    thyrotropin level of 0.04 µIU/mL | 0
    free thyroxine level of 1.64 ng/dL | 0
    normal free triiodothyronine level | 0
    peripheral blood leukocyte count of 11.58 × 109/L | 0
    78% neutrophils | 0
    erythrocyte sedimentation rate (ESR) of 95 mm/hour | 0
    ultrasound disclosed solid nodule with intranodular calcifications in the right thyroid lobe | 0
    outpatient diagnosis of subacute thyroiditis | 0
    treatment with cefixime 0.1 mg orally twice daily | -720
    treatment with ibuprofen 300 mg sustained-release capsules twice daily | -720
    poor treatment response | -720
    repeat thyroid function tests one month later | 0
    thyrotropin of 0.02 µIU/mL | 0
    free thyroxine of 35.0 pmol/L | 0
    free triiodothyronine of 5.3 pmol/L | 0
    thyroglobulin 78.93 ng/mL | 0
    thyroxine receptor antibody of 0.46 IU/L | 0
    peripheral blood leukocyte count of 16.87 × 109/L | 0
    peripheral blood leukocyte count increased to 22.46 × 109/L | 0
    86.9% neutrophils | 0
    ESR of 86 mm/hour | 0
    neuron-specific enolase level of 16.6 ng/mL | 0
    bone collagen CYFRA21-1 level of 11.16 ng/mL | 0
    ultrasound revealed diffuse thyroid disease suggestive of subacute thyroiditis | 0
    hypoechoic solid nodule with calcification in the right thyroid lobe | 0
    polyglandular lymphadenopathy with cortical thickening | 0
    medical history of Graves’ disease | -87600
    Graves’ disease complicated by hyperthyroidism | -87600
    adenomatoid thyroid nodules diagnosed via FNAC 2 years earlier | -17520
    chronic pharyngitis | -26280
    type II diabetes mellitus | -26280
    hypertension | -26280
    outmoded cerebral infarction | -26280
    pre-excitation syndrome | -26280
    denied radiation exposure | 0
    denied family history of thyroid diseases | 0
    denied family history of other malignancies | 0
    hospitalized | 0
    treated with oral prednisone acetate 10 mg twice daily | 0
    treated with rapid-acting insulin subcutaneously thrice daily after meals | 0
    treated with long-acting insulin subcutaneously at bedtime | 0
    treated with oral metformin 0.5 g thrice daily | 0
    treated with irbesartan 150 mg once daily | 0
    treated with nifedipine controlled-release tablets 30 mg once daily | 0
    treated with bisoprolol 5 mg once daily | 0
    treated with rosuvastatin 5 mg once nightly | 0
    treated with aspirin 100 mg once daily | 0
    prednisone tapered to 10 mg daily on day 16 | 384
    resolution of neck pain | 384
    insidious onset of dysphagia | 384
    choking cough | 384
    dyspnea | 384
    dysphonia | 384
    chest radiography disclosed right-sided tracheal deviation | 0
    computed tomography of the chest and neck revealed bilateral enlargement of the thyroid lobes and isthmus | 0
    heterogeneity and indistinct boundaries | 0
    tracheal stenosis | 0
    polyglandular lymphadenopathy involving bilateral supraclavicular nodes and perithyroid and carotid spaces | 0
    stroboscopic laryngoscopy disclosed limited movement of right vocal cord | 0
    limited movement of right arytenoid cartilage | 0
    normal left-sided function | 0
    both vocal cords closed | 0
    painless gastroscopy revealed stenotic esophageal entrance | 0
    partial thyroidectomy | 552
    tracheotomy performed under extracorporeal membrane oxygenation | 552
    postoperative pathological examination disclosed lesion with eggshell-calcified nodule | 552
    histopathologic evaluation revealed poorly differentiated malignant tumor | 552
    features of squamous cell carcinoma (SCC) | 552
    extensive necrosis with inflammatory reaction | 552
    invasion of adjacent striated muscle | 552
    invasion of vasculature | 552
    invasion of nerves | 552
    immunohistochemistry revealed galectin-3 (+) | 552
    cytokeratin 19 (CK19; +) | 552
    CD56 (−) | 552
    Ki-67 (70% +) | 552
    p53 (−) | 552
    TTF-1 (minority +) | 552
    TG (−) | 552
    calcitonin (−) | 552
    synuclein (−) | 552
    CGA (−) | 552
    Pax8 (+) | 552
    vimentin (scattered +) | 552
    final diagnosis of PSCCT | 552
    admitted to the intensive care unit postoperatively | 552
    tumor gradually metastasized to the lungs | 552
    metastasis to the face | 552
    metastasis to other anatomic sites | 552
    surgical site infection | 552
    multiple organ failures | 552
    wound infection progressed to sepsis | 552
    death | 552
    
    