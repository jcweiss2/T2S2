29 years old | 0
male | 0
admitted to the hospital | 0
hepatic transplantation | -4320
autoimmune hepatitis | -4320
minimal shortness of breath | 0
orthopnea | 0
loud superficial systodiastolic murmur | 0
palpable thrill | 0
edema | 0
ascites | 0
hypoalbuminemia | 0
thrombocytopenia | 0
hyperbilirubinemia | 0
ruptured aneurysm | 0
noncoronary sinus of valsalva | 0
turbulent flow | 0
aortic aneurysm | 0
left atrium | 0
mitral valve | 0
mild aortic regurgitation | 0
moderate mitral regurgitation | 0
continuous high-velocity jet | 0
cardiology and cardiovascular surgeon's council | 0
surgical operation recommended | 0
patient refused surgery | 0
hepatic transplant preparations delayed | 0
discharged | 168
elevated hepatic enzymes | 2160
ascites | 2160
diffuse edema | 2160
fever | 2160
infection parameters increased | 2160
complement values decreased | 2160
blood cultures | 2160
viridans group streptococcus | 2160
bedside portable echocardiography | 2160
gross vegetations | 2160
ampicillin initiated | 2160
gentamicin initiated | 2160
septic shock developed | 2160
multiple organ dysfunction syndrome | 2160
died | 2160