15 years old | 0
Saudi Arabian | 0
male | 0
presented to the emergency department | 0
vomiting | -72
headache | -72
hemoptysis | -72
shortness of breath | 0
referred from secondary care hospital | 0
intubated | 0
decreased oxygen saturation | 0
initial diagnosis of meningitis | 0
acute respiratory distress syndrome | 0
temperature 37.2°C | 0
heart rate 132 bpm | 0
blood pressure 135/95 mmHg | 0
crepitus at both upper regions of the chest | 0
no clinical abnormality in abdominal system | 0
no clinical abnormality in cardiovascular system | 0
laboratory findings of blood count not significant | 0
neck and chest contrast-enhanced CT revealed retropharyngeal abscess | 0
abscess extends to superior mediastinum | 0
abscess extends to posterior mediastinum | 0
marked mass effect on adjacent structures | 0
anterior displacement of pharynx | 0
anterior displacement of oesophagus | 0
anterior displacement of trachea | 0
conservative management | 0
no improvement | 24
surgical intervention | 24
pus drained from neck and mediastinal regions | 24
improvement on first post-operative day | 24
culture and sensitivity showed Ochrobactrum anthropi | 24
extubated | 48
discharged on eighth post-operative day | 192
remained well at 2-month follow-up | 1344
