43 years old | 0
    male | 0
    jaundice | -168
    nausea | -168
    vomiting | -168
    abdominal pain | -168
    flu-like syndrome | -168
    fever | -168
    chills | -168
    headache | -168
    myalgia | -168
    arthralgia | -168
    passing tea-colored urine | -168
    decreased urine output | -168
    asymptomatic chronic HBV infection | -96480
    treated as acute exacerbation of chronic HBV | -48
    transferred to our hospital | 0
    does not drink alcohol | 0
    alert | 0
    profound jaundice | 0
    abdominal upper quadrant tenderness | 0
    no hepatosplenomegaly | 0
    no ascites | 0
    normal neurological examination | 0
    acute kidney injury | 0
    creatinine 13.18 mg/dL | 0
    ureum 327 mg/dL | 0
    eGFR 4.06 mL/min/1.73m2 | 0
    elevated total bilirubin | 0
    indirect bilirubin 29.06 mg/dL | 0
    elevated liver transaminases | 0
    anemia | 0
    thrombocytopenia | 0
    hypoalbuminemia | 0
    positive bilirubin in urine | 0
    positive urobilinogen in urine | 0
    no hemoglobin detected in urine | 0
    polymerase chain reaction test negative for Covid-19 | 0
    positive HBsAg | 0
    positive IgM anti-HBc | 0
    positive anti-HBe | 0
    negative HBeAg | 0
    HBV-DNA quantification not performed | 0
    negative hepatitis C | 0
    negative hepatitis D | 0
    negative HIV | 0
    normal liver size | 0
    normal liver parenchyma | 0
    no splenomegaly | 0
    no ascites on ultrasound | 0
    severe liver fibrosis F3-F4 | 0
    median liver stiffness 14.9 kPa | 0
    treated with telbivudine | 0
    treated with cefoperazone | 0
    treated with furosemide | 0
    treated with ursodeoxycholic acid | 0
    supportive management | 0
    developed altered consciousness | 24
    metabolic acidosis pH 7.087 | 24
    HCO3− 3.0 mmol/L | 24
    oliguria <200 mL/24 hours | 24
    symptoms occurred 4 days after returning from Serui, Papua | -96
    rapid diagnostic test for malaria positive | 24
    peripheral blood smear showed intraerythrocytic P. falciparum | 24
    parasitemia 12.6% | 24
    diagnosis of severe malaria | 24
    intravenous artesunate | 24
    oral primaquine | 24
    transferred to intensive care unit | 24
    intubated | 24
    CRRT with CVVHDF initiated | 24
    initial downtrend in ureum | 24
    initial downtrend in creatinine | 24
    initial downtrend in bilirubin | 24
    initial downtrend in liver enzymes | 24
    improvement in eGFR | 24
    renal function continued to decline | 72
    liver injury deteriorated | 72
    developed pulmonary edema | 168
    developed septic shock | 168
    developed multiorgan dysfunction | 168
    died | 168
    negative malaria rapid test initially | 0
    positive malaria rapid test on day 2 | 24
    
    
    