69 years old|0
male|0
admitted to the ICU|0
pneumonia|0
severe sepsis|0
high doses of vasopressors|0
continuous hemodialysis|0
invasive ventilator support|0
remifentanil infusion|0
no long-acting opioids|0
weaned|336
decannulated|336
hyperactive delirium|336
confusion|336
paranoia|336
hallucinations|336
agitation|336
ICU delirium|336
no need for magnetic resonance imaging|336
non-pharmacological treatment|336
early mobility|336
sleep-wake cycle preservation|336
delirium persisted|336
prescribed 10 mg olanzapine orally|336
first prescription was 10 mg once daily|336
delirium worsened during the day|336
changed dosage to twice daily|336
fourth dose of olanzapine|0
awake|0
could recite his social security number|0
hypotensive|-30
blood pressure of 70/40 mmHg|-30
heart rate of 90 beats per min|-30
nonresponsive|-120
Glasgow coma scale score of 7|-120
pinpoint pupils|-120
maintained airway|-120
respiratory rate slightly elevated|-120
arterial blood gas showed normal pO2|-120
low pCO2|-120
blood sugar level slightly elevated|-120
norepinephrine infusion|-120
Glasgow coma scale score remained at 7|-120
ruled out hypoxia|-120
ruled out hypercapnia|-120
ruled out low blood sugar|-120
ruled out severe hypotension|-120
clinical suspicion of intoxication|-120
given 0.4 mg naloxone i.v.|-120
no effect|-135
given 0.5 mg flumazenil i.v.|?
