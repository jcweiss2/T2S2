64 years old| 0
man | 0
referred to the hospital | 0
cough | 0
chest X-ray findings with right pleural effusion | 0
right hilar mass | 0
significant facial edema | 0
chest computed tomography (CT) showed superior vena cava (SVC) syndrome | 0
transbronchial biopsy performed | -72
diagnosis of SCLC confirmed | -72
whole-body search indicated right hilar metastasis | 0
mediastinal metastasis | 0
right supraclavicular metastasis | 0
aortic metastasis | 0
superior mediastinal lymph node metastasis | 0
pleural effusion | 0
enhanced brain magnetic resonance imaging revealed no brain metastases | 0
no abnormal findings in the abdomen | 0
extensive SCLC diagnosed | 0
carboplatin and etoposide started as first-line treatment | 0
right pneumothorax observed | 96
chest tube drainage initiated | 96
ampicillin/sulbactam empirically administered | 144
fever developed | 144
right thoracic empyema developed | 144
febrile neutropenia (159·μL−1) developed | 192
treatment changed to meropenem with filgrastim | 192
pleural effusion culture showed meropenem-sensitive peptostreptococcus infection | 192
patient’s condition did not improve | 192
diarrhea appeared | 456
fecal culture results (CD toxin and CD antigen) negative | 456
diarrhea persisted | 456
fever persisted | 456
white blood cell counts surged | 504
bloody stools developed | 576
abdominal pain developed | 576
abdominal CT showed ascites | 576
intestinal retention | 576
intussusception in the ileocecal region | 576
abscess in the left hepatic lobe | 576
ileus suspected | 576
intestinal perforation suspected | 576
emergency surgery performed | 600
extensive necrosis of the colon found intraoperatively | 600
extensive colectomy performed | 600
colostomy performed | 600
septic shock occurred | 600
intensive care management performed | 600
meropenem changed to piperacillin/tazobactam, vancomycin, and micafungin | 600
fever continued | 600
systemic inflammation continued | 600
portal vein thrombosis developed | 672
anticoagulation therapy initiated | 672
Entamoeba histolytica trophozoites found in pathological specimens | 672
severe inflammatory cell infiltration of entire intestinal wall | 672
abscess formation with bleeding | 672
fibrin in some parts | 672
loss of continuity of the intestinal wall | 672
amoebic colitis diagnosed | 672
gastrointestinal perforation diagnosed | 672
liver abscess diagnosed | 672
portal vein thrombosis diagnosed | 672
no history of amoebiasis | 672
no sexual intercourse with homosexuals | 672
no contact with commercial sex workers | 672
no sexual intercourse with unspecified number of people | 672
traveled to the Philippines seven years prior | 672
traveled to West Coast of the United States | 672
traveled to Hawaii | 672
traveled to Shanghai 10 years prior | 672
metronidazole given orally | 792
patient’s general condition improved | 792
liver abscess size 36mm x 30mm | 792
percutaneous catheter drainage deemed difficult | 792
bacterial culture of right pleural effusion negative | 1176
chest tube removed | 1176
pleural effusion culture performed multiple times | 1176
no Entamoeba histolytica detected | 1176
chemotherapy for SCLC scheduled | 1176
paromomycin administered for 10 days | 1032
lower gastrointestinal endoscopy performed | 1464
lumen showed mild white mucus | 1464
residual redness observed | 1464
biopsy detected carcasses of amoebic trophozoites | 1464
patient’s general condition improved | 1464
liver abscess shrank on abdominal echo | 1464
amoebic dysentery cured | 1464
palliative radiotherapy performed | 1416
SVC syndrome exacerbated | 1416
second cycle of chemotherapy initiated | 2016
carboplatin dose reduced (AUC 5) | 2016
etoposide dose reduced (75 mg/m²) | 2016
four cycles of chemotherapy completed | 2016
partial response achieved | 2016
no recurrence of amoebic dysentery | 2016
