61 years old | 0
female | 0
diagnosed case of squamous cell carcinoma | 0
stage 1 oesophagus | 0
elective laparoscopic oesophagectomy | 0
gastric pull through operation | 0
preoperative assessment | -24
left ventricular function normal | -24
morphology normal | -24
transthorasic echocardiography | -24
anxiolysis | -24
benzodiazepines | -24
induction | 0
fentanyl-propofol | 0
intubated | 0
rocuronium | 0
isoflurane | 0
O2 nitrous | 0
rocuronium | 0
post-operative intensive care unit | 0
tachycardia | 10
hypotension | 10
patient ventilator asynchrony | 10
increased thoracic drain output | 10
bloody drain output | 10
low central venous pressure | 10
sinus tachycardia | 10
normal arterial blood gas analysis | 10
normal cardiac enzymes | 10
lower pCO2 levels | 10
crystalloid infusion | 10
colloid infusion | 10
vasopressor infusion | 10
noradrenaline | 10
analgesia | 10
sedation | 10
midazolam | 10
fentanyl | 10
re-exploration | 12
no obvious bleeding | 12
drains repositioned | 12
persistent need of vasopressor | 12
no fever | 12
no leukocytosis | 12
no increase in procalcitonin | 12
sterile blood cultures | 12
poor progression of r wave | 48
hypokinesia of the distal septum | 48
apical ballooning | 48
left ventricular peak mid cavity gradient | 48
ejection fraction 40% | 48
no mitral regurgitation | 48
no aortic regurgitation | 48
normal troponin I | 48
normal creatinine kinase | 48
high myoglobin | 48
high brain natriuretic peptide | 48
low molecular weight heparin | 48
aspirin | 48
statins | 48
dobutamine infusion | 60
T wave inversion | 60
normal troponin I | 60
normal CK level | 60
normal myoglobin | 60
high BNP | 60
left ventricular peak mid cavity gradient | 60
ejection fraction 30% | 60
surgical site sepsis | 120
death | 168
multi drug resistant abdominal sepsis | 168
combined cardiogenic and septic shock | 168