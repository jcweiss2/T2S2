48 years old | 0
male | 0
admitted to the hospital | 0
altered mental status | 0
found covered in urines and feces | -24
confused for the past day | -24
bed ridden during the last month | -720
cough | -720
diarrhea | -720
body temperature 35.8°C | 0
tachycardic | 0
tachypneic | 0
minimal accessory muscle use | 0
oxygen saturation 100% | 0
diminished breath sounds on the lung bases | 0
soft abdomen | 0
distended abdomen | 0
non-tender abdomen | 0
bilateral pitting edema | 0
acute hypoxemic respiratory failure | 1
tachypnea up to 40 breaths/min | 1
oxygen saturation 85% on room air | 1
intubated | 1
transferred to intensive care | 1
bilateral pleural effusions | 1
small pericardial effusion | 1
large heterogeneous splenomegaly | 1
ascites | 1
mesenteric and soft-tissue anasarca | 1
diffuse cerebral atrophy | 1
severe hyperferritinemia | 1
hyperferritinemia | 1
sepsis | 1
infections | 1
iron overload | 1
hepato-cellular disease | 1
kidney disease | 1
malignancy | 1
inflammatory/rheumatologic conditions | 1
blood cultures negative | 1
sputum cultures negative | 1
urine cultures negative | 1
HBsAg negative | 1
HBsAb negative | 1
hepatitis C antibody negative | 1
EBV PCR negative | 1
SARS-CoV-2 RNA PCR negative | 1
HIV 1,2 antigen/antibody test negative | 1
HTLV-1/2 antibodies negative | 1
CMV PCR ordered | 1
CMV PCR positive | 48
autoimmune workup negative | 1
diagnostic and therapeutic paracentesis | 48
diagnostic and therapeutic thoracentesis | 48
pleural fluid exudative | 48
pleural fluid lymphocytic | 48
cytology of pleural and ascitic fluids negative for malignant cells | 48
flow cytometry of pleural fluid showed T cell predominance | 48
T cell rearrangement study positive | 48
repeat chest CT suggestive of bilateral pneumonia | 48
bone marrow biopsy revealed histiocytes with hemophagocytic activity | 48
Interleukin 2 Receptor CD25 Soluble elevated | 48
diagnosis of HLH | 48
treated with fluids | 48
treated with vasopressors | 48
treated with broad-spectrum antibiotics | 48
renal replacement therapy initiated | 120
HLH-94 protocol initiated | 288
dexamethasone 20 mg daily | 288
renally adjusted etoposide 75 mg/m2 | 288
cardiac arrest | 298
pulseless electrical activity | 298
return of spontaneous circulation | 298
refractory shock | 304
died | 304
severe hyperkalemia | 304
hyperphosphatemia | 304
hypocalcemia | 304
hyperuricemia | 304
elevated blood urea nitrogen | 304
elevated creatinine | 304
TLS suspected | 304