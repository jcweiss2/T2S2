abdominal discomfort | -24
nausea | -24
vomiting | -24
no fever | -24
no vaginal discharge | -24
abdominal pain | -144
persistent nausea | -144
persistent vomiting | -144
tachycardia | -144
diffuse abdominal pain | -144
guarding on the right quadrants | -144
neutrophilia | -144
low prothrombinemia | -144
acute renal failure | -144
high procalcitonin | -144
high c-reactive protein | -144
moderate fluid in all quadrants | -144
good foetal vitality | -144
hypotension | -120
general abdominal guarding | -120
hyperlacticaemia | -120
hypokalaemia | -120
hyperglycaemia | -120
septic shock with an abdominal source | -120
emergency exploratory laparotomy | 0
generalised purulent peritonitis | 0
perforated acute appendicitis | 0
appendicectomy | 0
abdominal washing | 0
laparostomy | 0
admission to the Intensive Care Unit | 0
septic shock | 0
need for vasopressor therapy | 0
need for dialysis | 0
intravenous piperacillin-tazobactam antibiotherapy | 0
laparostomy revision | 48
marked bowel oedema | 48
bowel distention | 48
mild intraabdominal soiling | 48
further peritoneal lavage | 48
new laparostomy with progressive closure technique | 48
surgical revision | 96
abdominal cavity primary closure | 96
no need of prosthesis | 96
antibiotherapy adjustment | 144
piperacillin-tazobactam suspension | 144
amoxicillin with clavulanic acid initiation | 144
transfer to the obstetrics ward | 288
discharge home | 336
elective caesarean section | 1008
birth of a healthy child | 1008
ventral hernia | 936
obstetric follow-up | 936
good foetal viability | -24
good foetal vitality | -144 
daily evaluation by obstetrics physicians | 0 
good foetal viability | 0 
obstetric follow-up | 0 
no shortness of breath | -24 
denies chest pain | -24 
no neurological or other impairments | 936