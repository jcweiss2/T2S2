68 years old | 0
male | 0
obesity | 0
body mass index 34 kg/m2 | 0
admitted to the hospital | 0
acute respiratory failure | 0
fever | 0
respiratory rate 30/min | 0
pulse 80/min | 0
blood pressure 102/68 mmHg | 0
low oxygen saturation | 0
SpO2 85% on room air | 0
SARS-CoV-2 viral RNA negative | 0
Influenza A viral RNA negative | 0
Influenza B viral RNA negative | 0
pneumococcal urinary antigen negative | 0
hemocultures negative | 0
endotracheal intubation | 24
mechanical ventilation | 24
APACHE II score 18 | 24
chest CT scan | 24
bilateral infiltrates | 24
fibrosis | 24
coalescence | 24
SARS-CoV-2 anti-Spike IgG antibodies positive | 72
severe pneumonia due to COVID-19 | 72
ventilator-associated bacterial pneumonia | 216
Acinetobacter baumanii | 216
colistin therapy | 216
tigecycline therapy | 216
catheter-related A. baumanii bacteraemia | 408
colistin therapy | 408
tigecycline therapy | 408
tracheal aspirate positive for Pseudomonas putida | 888
blood culture positive for New Delhi metallo-β-lactamase 1 producing Enterobacter cloacae | 888
fosfomycin therapy | 888
gentamycin therapy | 888
tracheostomy | 1272
prone position | 1272
facial injuries | 1272
lower limbs injuries | 1272
sacral eschar grade III | 1272
bilateral nail hyperkeratosis lesions | 1272
fever | 1656
hemocultures | 1656
chest CT scan | 1656
Fusarium spp. | 1656
Fusarium verticillioides | 1656
antifungal therapy with amphotericin B | 1692
antifungal therapy with voriconazole | 1692
fungemia cleared | 1764
respiratory instability | 1920
sepsis | 1920
shock | 1920
death | 1920