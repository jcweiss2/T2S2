20 years old | 0
male | 0
Bahraini | 0
admitted to the hospital | 0
headache | -744
photosensitivity | -744
nausea | -744
left eye blurred vision | -744
generalised body fatigue | -744
limb weakness denied | -744
abnormal movements denied | -744
seizure denied | -744
loss of consciousness denied | -744
sensory manifestations denied | -744
MRI brain requested | 0
analgesia | 0
Multiplanar multisequential images taken | 0
postimage | 0
preimage contrast | 0
heterogeneously hyperintense lesion on T2-weighted images | 0
peripheral hypointensity | 0
optic chiasm compressed | 0
cavernous sinuses mildly compressed | 0
internal carotid artery blood flow spared | 0
T1 images with no contrast showed fluid level | 0
macroadenoma of pituitary gland | 0
haemorrhage | 0
mass effect on optic chiasm | 0
pituitary hormonal assessment | 0
loss of libido | 0
failure of erection | 0
polyuria | 0
polydipsia | 0
gynaecomastia denied | 0
change in body part size denied | 0
central hypogonadism | 0
central hypoadrenalism | 0
normal thyroid function | 0
mildly elevated level of prolactin | 0
hydrocortisone commenced | 0
cranial nerve abnormalities denied | 0
limb abnormalities denied | 0
gait abnormalities denied | 0
thyromegaly denied | 0
acromegaly denied | 0
chest X-ray normal | 0
trans-sphenoidal surgery | 744
incision done in the right nostril | 744
mucosa separated | 744
sphenoid sinus mucosa removed | 744
sellar floor identified | 744
sellar floor removed | 744
thick capsule of abscess incised | 744
yellowish pus drained | 744
cavity cleaned | 744
cavity irrigated with antibiotics and saline | 744
pus sent for Gram stain | 744
pus sent for culture | 744
pus sent for acid-fast bacilli stain | 744
pus sent for histopathological evaluation | 744
pituitary not removed | 744
histopathology showed inflammatory lesion | 744
histopathology showed no evidence of pituitary adenoma | 744
Gram stain showed few WBC | 744
culture sterile | 744
acid-fast bacilli stain negative | 744
metronidazole commenced | 744
ceftriaxone commenced | 744
vancomycin commenced | 744
antibiotics continued for 6 weeks | 744
patient doing well | 1488
symptoms improved | 1488
functional status normal | 1488
pituitary insufficiency continued | 1488
hydrocortisone continued | 1488
headaches denied | 1488
other symptoms denied | 1488
follow-up MRI | 1488
no enhancing residual abscess pockets | 1488
complete resolution | 1488