81 years old | 0
    female | 0
    multiple myeloma | 0
    dexamethasone | 0
    zoledronic acid | 0
    breast cancer | -87600
    lumpectomy | -87600
    radiation therapy | -87600
    hypertension | 0
    hypothyroidism | 0
    admitted | 0
    cough | -168
    runny nose | -168
    sore throat | -168
    denied fever | 0
    denied shortness of breath | 0
    denied chest pain | 0
    denied skin rashes | 0
    denied abdominal pain | 0
    denied diarrhea | 0
    tachypneic | 0
    no pharyngeal erythema | 0
    no tonsil exudates | 0
    no respiratory accessory muscle use | 0
    lungs clear | 0
    no skin rashes | 0
    white blood cell count 15.1 × 109/L | 0
    95% segmented neutrophils | 0
    bicarbonate 17 mmol/L | 0
    lactate 1.5 mmol/L | 0
    procalcitonin 0.28 ng/mL | 0
    chest radiograph no consolidations | 0
    computed tomography chest small airway disease | 0
    RSV positive | 0
    required 2 L oxygen | 0
    oxygen requirements increased | 48
    required high-flow oxygen | 48
    ribavirin started | 48
    transferred to ICU | 120
    intubated | 120
    respiratory distress | 120
    extubated | 216
    bilateral lower extremity weakness | 216
    absent lower extremity deep tendon reflexes | 216
    paresthesias of feet | 216
    weakness progressed | 216
    upper extremities involved | 240
    normal electrolytes | 240
    normal complete blood count | 240
    normal procalcitonin | 240
    alkaline phosphatase 62 U/L | 240
    alanine aminotransferase 22 U/L | 240
    aspartate aminotransferase 57 U/L | 240
    creatine kinase 198 U/L | 240
    attempted lumbar puncture | 240
    plasmapheresis initiated | 240
    five plasmapheresis treatments | 240
    minimal improvement quadriparesis | 240
    minimal improvement sensory nerve deficit | 240
    EMG low amplitude motor responses | 240
    axonal sensorimotor peripheral neuropathy | 240
    diminished extraocular movements | 264
    absent gag reflex | 264
    pupil asymmetry | 264
    intubated again | 264
    care withdrawn | 264
    