67 years old | 0
lady | 0
presented to the emergency department | 0
sudden onset right loin pain | 0
history of constant colicky pain | -12
radiating to the right loin | -12
vomiting | -12
denied urinary symptoms | 0
denied haematuria | 0
autoimmune liver cirrhosis | -131712
atrophic gastritis | -131712
Type 2 diabetes mellitus | -131712
hysterectomy | -43800
coronary artery bypass surgery | -43800
metformin | -131712
non-anaphylactic reactions to penicillin | -131712
non-anaphylactic reactions to intravenous contrast | -131712
pale | 0
temperature of 36.8 °C | 0
BP 141/72 | 0
pulse of 81 beats per minute | 0
right sided tenderness | 0
worse in the right upper quadrant | 0
worse in the right loin | 0
no crepitus | 0
anaemia | 0
Hb 9.8 g/dL | 0
impaired renal function | 0
urea 13.2 mmol/L | 0
creatinine 183 μmol/L | 0
HbA1c of 5.3% | 0
normal liver function tests | 0
prothrombin time elevated | 0
activated partial thromboplastin time elevated | 0
absence of neutrophil leucocytosis | 0
WCC 9 × 109/L | 0
trace of blood on urinalysis | 0
non-contrast CT of the kidneys, ureters and bladder arranged | 0
gas outlining the pelvicalyceal system of the right kidney | 0
perifascial gas tracking along the right ureter | 0
no discrete fluid collections | 0
no calculi | 0
blood cultures | 0
urine cultures | 0
intravenous antibiotics started | 0
intravenous fluids started | 0
radiological diagnosis of emphysematous pyelonephritis | 0
differential diagnoses | 0
blood specimens grew Escherichia coli | 0
urine specimens grew Escherichia coli | 0
sensitive to Meropenem | 0
addition of Metronidazole | 0
developed pyrexia | 0
developed tachycardia | 0
developed hypotension | 0
developed oliguria | 0
transferred to HDU | 0
C-reactive protein rise | 0
failed to mount inflammatory response | 0
leucocyte count of 6 g/dL | 0
platelet count dropped | 0
kidney function deteriorated | 0
creatinine rising to 258 μmmol/L | 0
falling platelet count | 0
severe sepsis | 0
end-organ failure | 0
emergency right nephroureterectomy | 0
open approach through right loin incision | 0
peritoneum opened | 0
free peritoneal fluid | 0
cirrhosis of the liver | 0
necrosis of the right renal pelvis | 0
necrosis of the ureter | 0
oedema in the retroperitoneum | 0
peri-ureteric gas | 0
no perinephric abscess | 0
no perinephric collection | 0
ureteric necrosis extended to lower third of right ureter | 0
right nephrectomy | 0
ligation of renal vessels | 0
kidney specimen with ureter placed in retroperitoneal space | 0
second incision made | 0
excision of diseased distal ureter | 0
removed en bloc with kidney | 0
retroperitoneal drain | 0
urethral catheter | 0
transferred to ICU | 0
histopathology confirmed microscopic parenchymal abscesses | 0
haemorrhagic infarction of ureteric mucosa | 0
serositis | 0
post-operative day 4 pyrexia | 96
CT abdomen and pelvis | 96
small bilateral pleural effusions | 96
normal post-operative changes | 96
no significant retroperitoneal collections | 96
smooth recovery | 312
IV antibiotics for 7 days | 168
discharged | 312
admission within 3 months of discharge | 1080
worsening renal function | 1080
managed conservatively | 1080
long term nephrology follow-up | 1080
