68 years old | 0
female | 0
admitted to the hospital | 0
incisional hernia | 0
history of repair of sigmoid perforation | -672
laparoscopic tension-free hernioplasty | 0
platelet count 224.1 × 10^9/L | 0
surgery was a success | 0
no excessive bleeding or hemorrhagic complications | 0
low platelet count 70.8 × 10^9/L | 96
shortness of breath | 96
chest tightness | 96
dizziness | 96
abdominal distension | 96
nausea | 96
low platelet count 36.9 × 10^9/L | 96
low white blood cell count 3.32 × 10^9/L | 96
culture from a purulent secretion revealed the growth of Escherichia coli | 96
serum endotoxin 54.51 pg/mL | 96
sepsis | 96
abdominal computed tomography scan showed extensive gas-fluid levels in the intestinal tract and intestinal wall swelling | 96
acute intestinal obstruction | 96
exploratory laparotomy | 120
intra-abdominal infections | 120
respiratory failure | 120
PaO2 51 mmHg | 120
PaCO2 45 mmHg | 120
transferred to the intensive care unit | 144
treated with fresh-frozen plasma | 144
treated with platelet transfusions | 144
treated with teicoplanin | 144
treated with ornidazole | 144
treated with imipenem | 144
treated with cilastatin sodium | 144
failed to respond to continuous platelet transfusions | 240
platelet count with EDTA 7.20 × 10^9/L | 240
platelet count with sodium citrate 136.00 × 10^9/L | 240
platelet clumps identified by microscopic examination | 240
EDTA-PTCP | 240
resolution of infection | 240
disappearance of EDTA-PTCP | 240