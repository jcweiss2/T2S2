81 years old| 0
    woman| 0
    hypertension| 0
    dyslipidemia| 0
    asthma| 0
    degenerative valve disease| 0
    presented to the emergency department| 0
    acute pre-cordial pain| 0
    dyspnea| 0
    nausea| 0
    vomiting| 0
    denied aspiration| 0
    hemodynamically stable| 0
    fever of 38.7 °C| 0
    signs of respiratory distress| 0
    hypoxemia| 0
    elevated inflammatory parameters| 0
    left pleural effusion| 0
    admitted| 0
    presumed diagnosis of aspiration pneumonia| 0
    began antibiotic treatment with amoxicillin| 0
    began antibiotic treatment with clavulanate acid| 0
    blood cultures were collected| 0
    elevation of the troponin level| 0
    peak 6.88 ng/mL| 0
    type 2 myocardial infarction| 0
    underwent transthoracic echocardiography| 0
    bad acoustic window| 0
    degenerative valve disease| 0
    moderate to severe aortic disease| 0
    important mitral valve calcification| 0
    moderate insufficiency| 0
    worsening of the dyspnea| 96
    worsening hypoxia| 96
    chest pain| 96
    chest computed tomography| 96
    excluded acute pulmonary embolism| 96
    extensive parenchymal consolidation of the left lung| 96
    antibiotic treatment altered to meropenem| 96
    combined with azithromycin| 96
    remained hypoxemic| 96
    worsening signs of respiratory distress| 96
    admitted to the intensive care unit| 96
    mechanically ventilated| 96
    new blood cultures were collected| 96
    developed circulatory shock| 96
    requiring noradrenalin| 96
    chest X-ray revealed bilateral infiltrates| 192
    underwent bronchofibroscopy| 192
    bronchial lavage| 192
    sputum collected for microbiology testing| 192
    blood cultures were negative| 192
    lavage cultures were negative| 192
    cycle of corticosteroids initiated| 192
    excessive post-infectious inflammatory process| 192
    interstitial lung disease| 192
    continued to worsen| 192
    febrile| 432
    chest X-ray revealed progressive lung infiltrates| 432
    steroids were suspended| 432
    TEE performed| 384
    confirmed important degenerative valve disease| 384
    severe aortic stenosis| 384
    P-MAIVF| 384
    important expansibility| 384
    solution of continuity| 384
    severe mitral regurgitation jet| 384
    mass in the tricuspid valve| 384
    probably due to infection| 384
    died| 480
    
    
    <|eot_id|>
    81 years old|0
    woman|0
    hypertension|0
    dyslipidemia|0
    asthma|0
    degenerative valve disease|0
    presented to the emergency department|0
    acute pre-cordial pain|0
    dyspnea|0
    nausea|0
    vomiting|0
    denied aspiration|0
    hemodynamically stable|0
    fever of 38.7 °C|0
    signs of respiratory distress|0
    hypoxemia|0
    elevated inflammatory parameters|0
    left pleural effusion|0
    admitted|0
    presumed diagnosis of aspiration pneumonia|0
    began antibiotic treatment with amoxicillin|0
    began antibiotic treatment with clavulanate acid|0
    blood cultures were collected|0
    elevation of the troponin level|0
    peak 6.88 ng/mL|0
    type 2 myocardial infarction|0
    underwent transthoracic echocardiography|0
    bad acoustic window|0
    degenerative valve disease|0
    moderate to severe aortic disease|0
    important mitral valve calcification|0
    moderate insufficiency|0
    worsening of the dyspnea|96
    worsening hypoxia|96
    chest pain|96
    chest computed tomography|96
    excluded acute pulmonary embolism|96
    extensive parenchymal consolidation of the left lung|96
    antibiotic treatment altered to meropenem|96
    combined with azithromycin|96
    remained hypoxemic|96
    worsening signs of respiratory distress|96
    admitted to the intensive care unit|96
    mechanically ventilated|96
    new blood cultures were collected|96
    developed circulatory shock|96
    requiring noradrenalin|96
    chest X-ray revealed bilateral infiltrates|192
    underwent bronchofibroscopy|192
    bronchial lavage|192
    sputum collected for microbiology testing|192
    blood cultures were negative|192
    lavage cultures were negative|192
    cycle of corticosteroids initiated|192
    excessive post-infectious inflammatory process|192
    interstitial lung disease|192
    continued to worsen|192
    febrile|432
    chest X-ray revealed progressive lung infiltrates|432
    steroids were suspended|432
    TEE performed|384
    confirmed important degenerative valve disease|384
    severe aortic stenosis|384
    P-MAIVF|384
    important expansibility|384
    solution of continuity|384
    severe mitral regurgitation jet|384
    mass in the tricuspid valve|384
    probably due to infection|384
    died|480