67 years old | 0
    male | 0
    admitted to the emergency department | 0
    left leg swelling | -168
    cactus plant injury | -168
    progressive left leg swelling | -48
    worsening erythema | -48
    pain | -48
    feeling generally unwell | -48
    blood pressure 71/41 mmHg | 0
    mean arterial pressure 48 mmHg | 0
    respiratory rate 36 breaths per minute | 0
    heart rate 125 beats per minute | 0
    sinus tachycardia | 0
    temperature 39°C | 0
    oxygen saturation 86% | 0
    admitted to the intensive care unit | 0
    pH 7.15 | 0
    PO2 84 mmHg | 0
    HCO3 15 mmol/L | 0
    lactate 7.6 mmol/L | 0
    sodium 134 mmol/L | 0
    urea 7.6 mmol/L | 0
    creatinine 173 μmol/L | 0
    eGFR 27 ml/min/1.73m² | 0
    white cell count 13.8 x10⁹/L | 0
    C-reactive protein 22 | 0
    hemoglobin 114 g/L | 0
    platelet 81 x10⁹/L | 0
    total bilirubin 99 μmol/L | 0
    ALT 61 U/L | 0
    AST 83 U/L | 0
    ALP 96 U/L | 0
    triple vasopressor support initiated | 0
    noradrenaline 20 mcg/min | 0
    adrenaline 20 mcg/min | 0
    vasopressin 0.04 units/min | 0
    piperacillin-tazobactam IV 4.5g | 0
    meropenem IV 2g | 0
    lincomycin IV 600mg | 0
    vancomycin IV 2g | 0
    emergency left lower limb fasciotomy | 0
    debridement | 0
    below knee amputation | 0
    LRINEC score 5 | 0
    left foot necrosis | 0
    below knee tissue necrosis | 0
    dishwasher fluid appearance | 0
    liquefied fat | 0
    unviable skin | 0
    unviable muscle | 0
    histopathology confirmed diagnosis | 0
    post-operative transfer to ICU | 24
    intubated | 24
    oliguria 10-14 ml/hour | 24
    pH 7.28 | 24
    lactate 4.7 mmol/L | 24
    sodium 130 mmol/L | 24
    creatinine 206 μmol/L | 24
    hemoglobin 89 g/L | 24
    platelet 105 x10⁹/L | 24
    white cell count 17 x10⁹/L | 24
    C-reactive protein 78 | 24
    INR 2.2 | 24
    APTT 150 sec | 24
    Group B Streptococcus pneumoniae isolated | 24
    ventilation sedation | 24
    propofol 170 mg/hr | 24
    fentanyl 40 mcg/hr | 24
    continuous renal replacement therapy initiated | 24
    noradrenaline 23 mcg/min | 24
    adrenaline 18 mcg/min | 24
    vasopressin 0.04 units/min | 24
    meropenem IV 2g TDS | 24
    lincomycin IV 600mg TDS | 24
    vancomycin IV 2g BD | 24
    IV immunoglobulin therapy 100g | 24
    surgical re-exploration | 24
    rapid atrial fibrillation | 48
    heart rate 110 bpm | 48
    oliguria 7@-25 ml/hour | 48
    pH 7.40 | 48
    lactate 3.9 mmol/L | 48
    sodium 131 mmol/L | 48
    creatinine 116 μmol/L | 48
    white cell count 26 x10⁹/L | 48
    C-reactive protein 105 | 48
    procalcitonin 21.18 μg/L | 48
    hemoglobin 83 g/L | 48
    platelet 63 x10⁹/L | 48
    INR 3.1 | 48
    fibrinogen 2.4 g/L | 48
    moderate left ventricular dysfunction | 48
    ejection fraction 40-45% | 48
    dilated atria | 48
    raised right atrial pressure | 48
    amiodarone loading dose 300mg | 48
    amiodarone maintenance dose 900mg | 48
    Oxiris filter applied | 48
    citrate anticoagulation circuit | 48
    sepsis-induced coagulopathy | 72
    surgical debridement | 72
    pH 7.31 | 72
    lactate 2.4 mmol/L | 72
    sodium 135 mmol/L | 72
    creatinine 79 μmol/L | 72
    white cell count 27 x10⁹/L | 72
    C-reactive protein 127 | 72
    hemoglobin 78 g/L | 72
    platelet 50 x10⁹/L | 72
    INR 2.0 | 72
    histopathology consistent with NF | 72
    wound culture growth of GBSPn | 72
    tissue culture growth of GBSPn | 72
    noradrenaline 20 mcg/min | 72
    adrenaline discontinued | 72
    vasopressin 2.4 units/min | 72
    refractory oliguria | 96
    furosemide IV 250mg | 96
    purpura over right forearm | 96
    weeping skin tears on right upper thigh | 96
    rapid atrial fibrillation HR 130 | 96
    pH 7.36 | 96
    lactate 1.5 mmol/L | 96
    sodium 130 mmol/L | 96
    creatinine 116 μmol/L | 96
    white cell count 33 x10⁹/L | 96
    C-reactive protein 103 | 96
    procalcitonin 15.37 μg/L | 96
    hemoglobin 91 g/L | 96
    platelet 53 x10⁹/L | 96
    INR 1.7 | 96
    bilirubin 131 μmol/L | 96
    AST 127 U/L | 96
    ALP 121 U/L | 96
    noradrenaline 20 mcg/min | 96
    vasopressin 2.4 units/min | 96
    amiodarone infusion | 96
    fulminant hepatic failure | 120
    encephalopathy | 120
    refractory oliguria 0@-5 ml/hour | 120
    pH 7.39 | 120
    lactate 1.2 mmol/L | 120
    sodium 134 mmol/L | 120
    creatinine 124 μmol/L | 120
    white cell count 39.5 x10⁹/L | 120
    C-reactive protein 74 | 120
    hemoglobin 116 g/L | 120
    platelet 49 x10⁹/L | 120
    INR 1.5 | 120
    bilirubin 139 μmol/L | 120
    AST 69 U/L | 120
    ALT 97 U/L | 120
    ALP 140 U/L | 120
    noradrenaline 20 mcg/min | 120
    vasopressin discontinued | 120
    ICU-acquired weakness | 144
    unarousable | 144
    no response to noxious stimuli | 144
    refractory oliguria 5 ml/hour | 144
    pH 7.44 | 144
    lactate 1.1 mmol/L | 144
    white cell count 43.5 x10⁹/L | 144
    C-reactive protein 109 | 144
    hemoglobin 90 g/L | 144
    platelet 57 x10⁹/L | 144
    INR 1.5 | 144
    bilirubin 150 μmol/L | 144
    AST 95 U/L | 144
    ALP 154 U/L | 144
    sedation discontinued | 144
    vasopressors discontinued | 144
    lincomycin discontinued | 144
    vancomycin discontinued | 144
    rifaximin 550mg BD | 144
    lactulose 20ml TDS | 144
    PRBC transfusion 2 units | 144
    jaundice | 168
    hypoactive delirium | 168
    RASS -5 | 168
    lateralizing signs to left | 168
    refractory oliguria | 168
    CT brain no acute pathology | 168
    acute calculous cholecystitis | 168
    pH 7.44 | 168
    lactate 1.1 mmol/L | 168
    white cell count 44.3 x10⁹/L | 168
    C-reactive protein 109 | 168
    hemoglobin 129 g/L | 168
    platelet 66 x10⁹/L | 168
    INR 1.3 | 168
    bilirubin 235 μmol/L | 168
    AST 75 U/L | 168
    ALP 175 U/L | 168
    conjugated bilirubin 142 μmol/L | 168
    meropenem continued | 168
    anuria | 192
    hypotensive BP 71/33 mmHg | 192
    MAP 51 mmHg | 192
    febrile 39°C | 192
    rapid atrial fibrillation HR 160 | 192
    troponin 616 | 192
    ammonia 158 μmol/L | 192
    bilirubin 352 μmol/L | 192
    AST 100 U/L | 192
    ALP 299 U/L | 192
    furosemide IV 250mg | 192
    acetazolamide IV 500mg | 192
    noradrenaline 2.5 mcg/min | 192
    lincomycin IV 600mg TDS | 192
    digoxin IV 500mcg | 192
    metoprolol IV 15mg | 192
    palliative care pathway | 192
    deceased | 192
