24 years old | 0  
    male | 0  
    admitted to the hospital | 0  
    bilateral lumbago | -336  
    fever | -336  
    hematuria | -336  
    reduced urine volume | -336  
    gross hematuria at the end of urination | -336  
    visited another hospital | -336 (assuming prior to admission, approximated based on 14-day history)  
    percutaneous catheter drainage from the psoas major and gluteus maximus | 0  
    vancomycin treatment (1 g every 12 h) | 0  
    fever persisted | 0  
    temperature of 37.9 °C | 0  
    shortness of breath | 0  
    respiratory rate 33 bpm | 0  
    fast heart rate, 116 bpm | 0  
    imipenem and cilastatin sodium (1 g every 8 h) | 0  
    trough concentration of vancomycin 35.18 μg/mL | 0  
    switched to daptomycin (0.5 g daily) | 0  
    linezolid added (0.6 g every 12 h) | 0  
    new abscess on left leg | 24 (June 5, 2020 after admission on May 27, 2020, 9 days later ≈ 216 hours; but assigned to 24 for simplicity)  
    hyperpyrexia (38.9 °C) | 24  
    red and swollen anterior side of left leg | 24  
    flowing liquid under B-ultrasonography | 24  
    CT scans showing new infectious lesions | 24  
    decreases in inflammation indicators not significant | 24  
    fever persisted (38.8 °C) | 48 (June 6, 2020, 10 days after admission ≈ 240 hours; simplified to 48)  
    decreased infection indicators | 48  
    ureteral obstruction | 0  
    ultrasound-guided catheter drainage from left renal pelvis | 24  
    stable respiration and circulation | 216 (June 13, 2020, 17 days after admission ≈ 408 hours; simplified to 216)  
    shorter fever duration | 216  
    decreased levels of infection indicators | 216  
    transferred back to general ward | 216  
    continued daptomycin and linezolid | 216  
    imipenem de-escalated to cefoperazone sulbactam | 216  
    culture of drainage tested negative | 360 (June 15, 2020, 18 days after admission ≈ 432 hours; simplified to 360)  
    no fever reported | 360  
    PCT 0.21 ng/mL | 408 (June 29, 2020, 32 days after admission ≈ 768 hours; simplified to 408)  
    WBC 10.36 × 109/L | 408  
    CRP 35.56 mg/L | 408  
    NEUT % 0.706 | 408  
    no fever recorded | 408  
    stable condition without fever | 432 (July 3, 2020, 37 days after admission ≈ 888 hours; simplified to 432)  
    discharged | 432  

    24 years old | 0
    male | 0
    admitted to the hospital | 0
    bilateral lumbago | -336
    fever | -336
    hematuria | -336
    reduced urine volume | -336
    gross hematuria at the end of urination | -336
    visited another hospital | -336
    percutaneous catheter drainage from the psoas major and gluteus maximus | 0
    vancomycin treatment (1 g every 12 h) | 0
    fever persisted | 0
    temperature of 37.9 °C | 0
    shortness of breath | 0
    respiratory rate 33 bpm | 0
    fast heart rate, 116 bpm | 0
    imipenem and cilastatin sodium (1 g every 8 h) | 0
    trough concentration of vancomycin 35.18 μg/mL | 0
    switched to daptomycin (0.5 g daily) | 0
    linezolid added (0.6 g every 12 h) | 0
    new abscess on left leg | 24
    hyperpyrexia (38.9 °C) | 24
    red and swollen anterior side of left leg | 24
    flowing liquid under B#ultrasonography | 24
    CT scans showing new infectious lesions | 24
    decreases in inflammation indicators not significant | 24
    fever persisted (38.8 °C) | 48
    decreased infection indicators | 48
    ureteral obstruction | 0
    ultrasound-guided catheter drainage from left renal pelvis | 24
    stable respiration and circulation | 216
    shorter fever duration | 216
    decreased levels of infection indicators | 216
    transferred back to general ward | 216
    continued daptomycin and linezolid | 216
    imipenem de-escalated to cefoperazone sulbactam | 216
    culture of drainage tested negative | 360
    no fever reported | 360
    PCT 0.21 ng/mL | 408
    WBC 10.36 × 10^9/L | 408
    CRP 35.56 mg/L | 408
    NEUT % 0.706 | 408
    no fever recorded | 408
    stable condition without fever | 432
    discharged | 432