18 years old | 0
male | 0
attended a health center | 0
fatigue | -24
anosmia | -24
dyspnea | -24
SpO2 levels 55% | -24
SpO2 levels 75% | -24
hospitalized | -24
chest radiography | -24
bilateral lung infiltrates | -24
RT-PCR swab tested positive for SARS-CoV-2 infection | -24
admitted in a COVID-19 infirmary unit | -24
non-invasive ventilation support | -24
intubation and invasive mechanical ventilation | -24
ventral decubitus positioning | -24
Escherichia coli | -48
methicillin-sensitive Staphylococcus aureus | -48
amoxicillin | -48
blood culture revealed methicillin-resistant Staphylococcus aureus | -48
dismissed | -48
clinical improvement | -48
extubated | -48
discharged | -48
attended the emergency department | -336
retrosternal thoracalgia | -336
irradiating to the left upper limb | -336
soft tissue swelling of the shoulder and arm | -336
fever | -336
increased levels of C-reactive protein | -336
hemoculture and urine culture proved negative | -336
chest radiograph and thoracic CT | -336
typical changes compatible with sequelae of Covid-19 pneumonia | -336
admitted for further investigation and treatment planning | -336
gentamicin | -336
prescribed and administered | -336
thoracic CT with intravenous contrast administration | -345
scapulohumeral synovitis | -345
multiple intra-muscular collections | -345
glenohumeral joint | -345
scapulohumeral synovitis and less pronounced joint fluid | -345
bilateral shoulder magnetic resonance imaging (MRI) with intravenous contrast administration | -396
infraspinatus fossa and subscapular fossa collections | -396
capsular thickening and increased signal intensity post-gadolinium administration | -396
septic arthritis and rotator cuff collections | -396
myonecrosis | -396
aspiration of the infraspinatus fossa collection | -408
seropurulent fluid | -408
8,5 Fr drainage catheter | -409
removed | -409
evaluation of the aspirate | -409
direct and culture tests for Mycobacterium tuberculosis, anaerobic and aerobic bacteria | -409
negative | -409
improvement of left shoulder range of motion | -408
physical rehabilitation exercises | -408
transferred to another hospital | -408
continue physical therapy and rehabilitation exercises | -408
prolonged immobilization | -24
mechanical ventilation | -24
muscle atrophy | -24
heterotopic ossification around the shoulder | -24
delirium | -24
lung damage | -24
muscle weakness | -24
rhabdomyolysis | -336
myalgia | -336
fatigue | -336
pigmenturia | -336
acute renal failure | -336
imaging findings | -336
enlargement of the affected muscles | -336
MRI | -408
hyperintense signal on fluid-sensitive sequences | -408
heterogeneous enhancement following intravenous contrast administration | -408
rim enhancement | -408
septic arthritis | -336
arthralgia | -336
muscle pain | -24
fatigue | -24
arthropathy | -24
arthropathy excluded | -336
antibiotic regimen | -336
unknown cause of bilateral shoulder arthritis | -336
presumed of septic nature | -336