83 years old | 0
male | 0
admitted to the emergency facility | 0
dislodgment of gastrostomy feeding tube | -24
gastrostomy | -648
swallowing disorder | -648
acute ischemic stroke | -648
stoma was stenotic | 0
dilation of stoma | 0
new tube inserted | 0
abdominal pain | 1
vomiting | 1
diet administration | 1
returned to the hospital | 36
physical examination | 36
ill-looking patient | 36
dehydrated | 36
hypotension | 36
tachycardia | 36
abdomen was distended | 36
diffusely tender | 36
abdominal computed tomography (CT) | 36
infusion of iodine contrast medium | 36
cavity formed by peritoneal blockade | 36
exploratory laparotomy | 36
surgical findings | 36
lumpy liquid in the peritoneal cavity | 36
peritoneal adhesions | 36
false path | 36
blockade purulent collection | 36
another gastrostomy | 36
stomach sutured to the abdominal wall | 36
thorough lavage of the peritoneal cavity | 36
abdomen was drained | 36
referred to the intensive care unit | 36
evisceration | 37
re-operation | 37
multiple organ failure | 43
death | 43
periostomal infection | -648
stomal leakage | -648
tube dislodgment | -24
severe wound infection | 36
septicemia | 36
dehiscence | 37
aspiration | 36
peritonitis | 36
gastrointestinal perforation | 36
bleeding | 36
skin ulceration | -648
superficial abscesses | -648
retrograde jejunoduodenogastric intussusception | -648