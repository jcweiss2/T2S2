42 years old | 0
    man | 0
    presented to our center | 0
    high-grade fever | -1008
    chills | -1008
    productive cough since six weeks | -1008
    weight loss (6 kg over four weeks) | -672
    diarrhea since two weeks | -336
    chest radiograph (CXR) showed right middle zone consolidation | -4320
    sputum culture grew Klebsiella pneumoniae | -4320
    antibiotics were started (levofloxacin, amikacin, metronidazole, fluconazole) | -4320
    empiric anti-tuberculosis therapy (ATT) was started | -4320
    referred to our hospital | -4320
    asymptomatic until 5 years ago | -43440
    recurrent upper respiratory tract infections (RTIs) since 2005 | -43440
    pneumonia (2006) | -43440
    treated for pulmonary tuberculosis twice (2005, 2007) | -43440
    monthly episodes of watery diarrhea since 2007 | -43440
    childhood and family history were insignificant | 0
    examination revealed fever | 0
    tachycardia | 0
    tachypnea (respiratory rate 36/min) | 0
    blood pressure of 110/60 | 0
    bilateral crepitations on chest auscultation | 0
    PaO2 was 58 mm Hg on arterial blood gas analysis | 0
    admitted to the intensive care unit (ICU) | 0
    CXR showed right middle and lower zone consolidation | 0
    non-resolving pneumonia (NRP) was diagnosed | 0
    meropenem and levofloxacin were started | 0
    ATT discontinued | 0
    endotracheal intubation was soon required | 0
    CXR showed bilateral alveolar shadows | 120
    PaO2/FiO2 of 59/1 (<200) | 120
    ventilation with ARDS protocol was started | 120
    noradrenaline was given at ceiling doses | 120
    antibiotics were changed (targocid, colistin) | 120
    empiric amphotericin-B was added | 120
    trimethoprim-cotrimoxazole prophylaxis was started | 120
    underlying primary immune deficiency (PID), a CVID, was suspected | 168
    intravenous immunoglobulin (IVIG) was given (2 g/kg on 21/9/09) | 168
    hypogammaglobulinemia | 168
    became afebrile for the first time in eight weeks | 192
    FiO2 requirements reduced (35% by 6/10/09) | 192
    tracheostomy was done (30/10/09) | 1296
    subsequent decannulation (26/10/09) | 1248
    CXR showed clearing of alveolar shadows | 1248
    residual bronchiectasis | 1248
    ambulatory on discharge | 1248
    follows up (irregularly, due to cost constraints) for replacement IVIG and chest physiotherapy | 1248
    serum immunoglobulin level measurement | 0
    low CD4 T lymphocyte counts | 0
    HIV infection ruled out | 0
    recurrent RTIs and diarrhea, beginning 5 years prior to presentation | -43440
    infection with Klebsiella pneumoniae and Pseudomonas aeruginosa | 0
    IVIG commenced (2 g/kg loading dose, over 5 days) | 168
    significant improvement followed within 72 hours | 192
    repeat IgG levels after 8 and 12 weeks of loading dose | 1248
    replacement doses (0.4 g/kg) given | 1248
    confirming the diagnosis of a CVID | 1248
    recurrent RTIs | -43440
    chronic sinusitis | -43440
    lung fibrosis | -43440
    bronchiectasis (12.2%) | -43440
    granulomatous interstitial lung disease | -43440
    autoimmune phenomena | -43440
    systemic lymphocytic infiltration | -43440
    antibody deficiency | -43440
    encapsulated bacteria infections | -43440
    IVIG replacement | 1248
    hypogammaglobulinemia treatment | 1248
    monthly dose of 0.4 g/kg | 1248
    maintenance of serum IgG trough level >0.8 g/l | 1248
    antibody failure precludes vaccine use | 0
    late-onset common immune deficiency category | 1248
    NRP with Gram-negative sepsis | 0
    ICU mortality of severe pneumonias was 36.8% | 0
    PIDs may be missed as a cause of NRPs | 0
    malnutrition | 0
    HIV infection | 0
    tuberculosis | 0
    inappropriate use of antibiotics | 0
    CVIDs are the most common PID | 0
    pneumonia deteriorated despite appropriate antibiotics, mechanical ventilation, and inotropes | 0
    CVIDs are an important cause of severe pneumonia even in adults | 0
    correct diagnosis and prompt treatment of underlying CVIDs can reduce mortality | 0
    source of support: Nil | 0
    conflict of interest: None declared | 0
    