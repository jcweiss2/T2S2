34 years old | 0
male | 0
transferred to intensive care unit | 0
pulmonary hemorrhage | 0
septic shock | 0
admitted to local hospital | -24
acute dyspnea | -24
hemoptysis | -24
fatigue | -168
back pain | -168
abdominal pain | -168
nausea | -168
vomiting | -168
temperature 35.9°C | -24
systolic blood pressure 70 mmHg | -24
heart rate 100 beats per minute | -24
respiratory rate 19 breaths per minute | -24
oxygen saturation 60% | -24
jaundice | -24
hemoptysis persisted | -24
abdominal pain over right upper quadrant | -24
chest auscultation revealed ubiquitous coarse crackles | -24
chest X-ray showed bilateral patchy infiltrates | -24
mild normochromic normocytic anemia | -24
hemoglobin 13.0 g/dL | -24
bilirubin 8.45 mg/dL | -24
severe thrombocytopenia 20×10^9/L | -24
acute renal failure | -24
creatinine level 4.9 mg/dL | -24
leukocytosis 31×10^9/L | -24
elevated C-reactive protein | -24
elevated procalcitonin levels | -24
diagnosis of community acquired pneumonia | -24
diagnosis of sepsis | -24
transferred to intensive care unit (primary hospital) | -24
blood cultures obtained | -24
empiric antimicrobial therapy with piperacillin/tazobactam | -24
empiric antimicrobial therapy with ciprofloxacin | -24
hypoxia aggravated | -16
non-invasive ventilation | -16
endotracheal intubation | -16
insufficient oxygenation despite mechanical ventilation | -16
ECMO therapy initiated | -16
ECMO team implanted venovenous ECMO | -16
transferred to tertiary referral hospital | 0
blood gases showed metabolic and respiratory acidosis | 0
blood gases showed hypoxemia | 0
CT-scan showed ARDS | 0
bronchoscopy revealed diffuse alveolar hemorrhage | 0
hemoptysis persisted | 0
intravascular hemolysis | 0
hemoglobin drop from 13.0 to 5.9 g/dL | 0
reduced haptoglobin | 0
increased lactate dehydrogenase | 0
coagulation compromised | 0
fibrinogen below 30 mg/dL | 0
transfusion of 10 packed red blood cells | 0
transfusion of 12 g fibrinogen | 0
hemoglobin stabilized at 7.0 g/dL | 0
urinalysis showed muddy-brown casts | 0
urinalysis showed acanthocytes | 0
hyperkalemia | 0
continuous venovenous renal replacement therapy | 0
citrate anticoagulation | 0
gastrointestinal symptoms prior to admission | 0
plasmapheresis initiated | 0
suspected hemolytic uremic syndrome | 0
volume therapy 13 L within 16 h | 0
sodium bicarbonate 2250 mL | 0
conventional therapy failed | 0
rescue therapy with extracorporeal cytokine absorbent filter | 0
prednisolone 1000 mg administered | 0
died in fulminant multi-organ failure | 17
fibrin monomers negative | 17
anti-glomerular basement antibodies negative | 17
anti-nuclear antibodies negative | 17
anti-neutrophil cytoplasmic antibodies negative | 17
peripheral blood smear detected 6–8% schistocytes | 17
ADAMTS-13 activity 35% | 17
LipL32-PCR positive for Leptospira interrogans | 24
blood cultures sterile | 24
urine samples sterile | 24
bronchoalveolar lavage samples sterile | 24
transmitted by pet rat | 0
purchased pet rat 4 weeks before admission | -672
Leptospira interrogans detected in rat kidney | 0
Plasmapheresis | 0
cortisone therapy | 0
beta-lactam antimicrobial therapy | 0
extracorporeal cytokine absorbent therapy | 0
no improvement in outcome | 17
diagnosis of leptospirosis | 24
death occurred 29 hours after initial presentation | 29
