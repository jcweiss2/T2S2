73 years old | 0
male | 0
admitted to the emergency department | 0
previous bioprosthetic aortic valve replacement | -131400
B-cell lymphoma | 0
active B-cell lymphoma | 0
newly diagnosed B-cell lymphoma | 0
receiving chemotherapy | 0
cardiogenic shock | 0
prosthetic heart valve failure | 0
acute aortic regurgitation | 0
infective endocarditis | 0
negative blood cultures | -72
transfemoral valve-in-valve TAVR | 168
balloon-expandable Edwards Sapien 3 heart valve | 168
general anesthesia | 168
excellent immediate procedural result | 168
full recovery | 168
prolonged suppressive antibiotic therapy | 168
septicemia | 0
embolic stroke | 0
systemic embolization | 0
septic shock | 0
mobile vegetations | 0
floating vegetations | 0
abscess | 0
fistula formation | 0
leaflet destruction | 0
cusp destruction | 0
prosthetic heart valve endocarditis | 0
inconclusive imaging | 0
transthoracic echocardiography | 0
transesophageal echocardiography | 0
multidetector-row CT | 0
FDG PET/CT | 0
relapsing infection | 0
recurrent endocarditis | 0
multiorgan failure | 0
cerebral embolism | 0
bridge to surgical repair | 0
parenteral antibiotic therapy | 0
incomplete device extraction | 0
device extraction | 0
sterilized valvular structures | 0
sterilized perivalvular tissues | 0
cardiac radionuclide imaging | 0
embolic stroke |;0
