72 years old | 0
male | 0
hypertension | 0
stage 3 chronic kidney disease | 0
abdominal discomfort | -672
constipation | -672
worsening oral intake | -672
somnolent | 0
diffuse abdominal pain | 0
afebrile | 0
tachypneic | 0
tachycardic | 0
white blood cell count 27.7 | 0
potassium 7.0 mmol/L | 0
metabolic acidosis CO2 11mmol/L | 0
AKI | 0
BUN 174 mg/dL | 0
creatinine 15.4 mg/dL | 0
microscopic urinalysis positive for >150 RBC and WBC per high power field | 0
few bacteria | 0
CT of the abdomen and pelvis | 0
multiple fluid collections | 0
gas throughout the abdomen | 0
pockets adjacent to the superior and posterior walls of the urinary bladder | 0
fleet enema | -72
surgical consultation | 0
suspected intestinal rupture | 0
interventional radiology guided fluid drainage | 0
broad spectrum antibiotics | 0
emergent hemodialysis | 0
ascitic analysis | 72
fluid Cr of 7 mg/dL | 72
bacterial culture positive for E. coli | 72
CT cystogram | 72
bladder rupture | 72
urinary bladder leakage | 72
intraperitoneal spillage of contrast | 72
open repair of the urinary bladder | 96
exploratory laparotomy | 96
two intestinal abscesses | 96
inflammation of the distal sigmoid | 96
inflammation of the appendix | 96
inflammation of the viscera | 96
drainage of abscesses | 96
prophylactic appendectomy | 96
diverting sigmoid colostomy | 96
vasodilatory shock | 96
vasopressors | 96
antimicrobial therapy | 96
renal recovery | 240
discharged | 240
sepsis secondary to UTI | 480
intra-abdominal fluid collection | 480
IV antibiotics | 480
discharged with a foley catheter | 480