60 years old | 0
male | 0
admitted to the hospital | 0
diabetes mellitus | 0
hypertension |A0
transurethral resection of the prostate | 0
refractory urine retention | 0
no loin pain | 0
no fever | 0
no rigors | 0
no previous surgery | 0
no renal angle tenderness | 0
benign digital rectal examination | 0
persistent pus cells (14/HPF) | 0
positive pansensitive Escherichia coli | 0
antibiotics (levofloxacin) | 0
urethral catheter exchange | 0
urinary tract ultrasound showed enlarged prostate of 46 gm | 0
transurethral resection of the prostate under antibiotic coverage (piperacillin/tazobactam) | 0
postoperative recurrent high-grade fever | 24
left loin pain | 24
elevated septic parameters | 24
urine culture positive for Candida albicans | 24
blood culture positive for Candida albicans | 24
intravenous fluconazole | 24
no response to fluconazole | 24
CT urography showed left hydronephrosis | 48
CT urography showed filling defect in left renal pelvis | 48
suspected renal fungal ball | 48
left percutaneous nephrostomy | 72
nephrostogram showed filling defects in renal pelvis | 72
whitish debris in nephrostomy urine | 72
whitish debris in urethral catheter urine | 72
cultures from nephrostomy positive for Candida albicans | 72
cultures from urethral catheter positive for Candida albicans | 72
cultures from blood positive for Candida albicans | 72
fever did not subside with intravenous fluconazole | 72
treatment changed to anidulafungin 100 mg once daily | 72
patient improved | 168
repeated blood culture negative | 168
urine from bladder positive for candida | 168
urine from nephrostomy positive for candida | 168
instillation of fluconazole through nephrostomy | 168
urine culture from nephrostomy tube showed no growth | 264
midstream urine showed mixed growth with some candida | 264
follow-up renal ultrasound showed normal left kidney | 264
nephrostomy tube removed | 336
urine culture one week later showed no candida growth | 336
Candida albicans infection | 0
fungal ball | 0
sepsis | 0
percutaneous nephrostomy | 72
intravenous antifungal agent | 72
fluconazole instillation | 168
no enhancement on CT urography | 48
contrast outlining the lesion with no attachment to renal pelvis | 48
diabetes mellitus as risk factor | 0
indwelling urethral catheter as risk factor | 0
use of antibiotics as risk factor | 0
community-acquired infection before hospitalization | 0
Candida albicans most common species | 0
urinary drainage devices as risk factor | 0
candiduria treatment recommended | 0
fluconazole and amphotericin B common | 0
echinocandins limited use | 0
relieve obstruction required | 72
local antifungal irrigation | 168
amphotericin B nephrotoxicity | 0
fluconazole instillation success | 168
treatment success indicators | 264
renal fungal ball rare | 0
management options include intravenous agents and percutaneous nephrostomy | 72
antifungal irrigation via nephrostomy | 168
conflicts of interest none | 0
