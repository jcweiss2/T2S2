71 years old | 0
woman | 0
chronic obstructive pulmonary disease | 0
atrial fibrillation | 0
bladder cancer | 0
type 2 insulin-dependent diabetes mellitus | 0
urinary tract infection | -168
surgery to resect bladder tumor | -672
UTI progressed to sepsis | -168
required transfer to intensive care unit | 0
home dose of 30 units per day of glargine insulin | -24
insulin sliding scale | -24
blood glucose became unresponsive to home insulin | 0
developed hyperosmolar hyperglycemic state |1
normal anion gap | 0
normal pH | 0
sodium level was normal | 0
increasing glargine dose | 24
blood glucose remained uncontrolled | 24
aspart boluses | 24
NPH boluses | 24
transitioned to regular insulin drip | 48
insulin drip lost efficacy | 72
insulin drip titrated up to maximum dose of 1620 units | 96
blood glucose remained above 400mg/dL | 96
test for insulin autoantibodies | 120
insulin autoantibodies negative | 120
theories for lack of insulin efficacy | 144
