76 years old | 0
female | 0
Caucasian | 0
admitted to hospital | 0
hypertension | -8760
dyslipidaemia | -8760
palpitations | -336
orthopnoea | -336
shortness of breath | -336
New York Heart Association functional class III–IV | -336
atrial fibrillation | 0
left bundle branch block | 0
decompensated heart failure | 0
pulmonary oedema | 0
bilateral pleural effusions | 0
intubated | 24
cardiac catheterization | 24
no flow-limiting stenoses | 24
right coronary artery emptying into pulmonary artery | 24
transthoracic echocardiogram | 24
severely reduced RV systolic function | 24
severe right atrial dilatation | 24
severe tricuspid regurgitation | 24
positive cultures for Streptococcus bovis | 48
intermittent haemodialysis | 168
transoesophageal echocardiogram | 216
dilated and tortuous left main coronary artery | 216
dilated and tortuous vessel draining into pulmonary artery | 216
anomalous right coronary artery from pulmonary artery | 216
turned down for surgical intervention | 216
transferred to hospice care | 960
deceased | 1800
uncontrolled atrial fibrillation | 0
left bundle branch block | 0
clinical evidence of decompensated heart failure | 0
chest X-ray confirming evidence of pulmonary oedema | 0
bilateral pleural effusions | 0
intravenous diuresis | 0
rate control | 0
increased WBC count | 8
eosinophilia | 8
systemic involvement | 8
fever | 8
diaphoretic | 8
tachycardic | 8
hypotensive | 8
high-sensitivity troponin increased | 8
serum lactate increased | 8
anuric acute kidney injury | 8
dual antiplatelet therapy | 8
vasopressors | 8
point-of-care ultrasound | 8
biventricular systolic dysfunction | 8
plethoric non-collapsible inferior vena cava | 8
diastolic flattening of the interventricular septum | 8
volume overload of the right ventricle | 8
ad hoc right heart catheterization | 24
haemodynamic assessment | 24
oximetry run | 24
no intra-cardiac left-to-right shunt | 24
pulmonary artery angiography | 24
no pulmonary embolus | 24
no fistula involving the RVOT | 24
pulmonary vascular resistance | 24
systemic vascular resistance | 24
RV angiogram | 24
significant tricuspid regurgitation | 24
dilated and severely dysfunctional right ventricle | 24
elevated cardiac index | 24
sepsis | 24
empiric antibiotics | 24
extubated | 240
transferred to cardiology ward | 240
intermittent haemodialysis | 240
dependent on intermittent haemodialysis | 240
no expected renal recovery | 240
potential therapeutic options for ARCAPA | 240
discussed at interdisciplinary heart team rounds | 240
not a surgical candidate | 240
pursue comfort measures | 240
cessation of dialysis | 240
transferred to hospice | 960
passed away | 1800