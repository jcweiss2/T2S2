67 years old | 0
male | 0
hypertension | -7200
benign prostatic hyperplasia | -7200
childhood asthma | -7200
admitted to the hospital | 0
abdominal pain | -672
bloating | -672
decreased oral intake | -672
shortness of breath | -672
fatigue | -672
no bowel movement | -72
denies fever | -672
denies chills | -672
denies cough | -672
denies trauma | -672
denies weight loss | -672
denies nausea | -672
denies vomiting | -672
denies diarrhea | -672
denies sick contacts | -672
denies recent travel | -672
denies hematuria | -672
denies hematochezia | -672
retired office manager | -7200
former smoker | -7200
drinking two to three beers every day | -7200
migrant from Cuba | -7200
living in the USA | -7200
finasteride | -7200
omeprazole | -7200
tamsulosin | -7200
afebrile | 0
blood pressure 102/47 mm Hg | 0
heart rate 149 beats per minute | 0
saturating well on room air | 0
bilateral decreased breath sounds | 0
wheezing at bases | 0
tachycardia | 0
irregularly irregular pulse | 0
trace bilateral pedal edema | 0
soft, mildly distended abdomen | 0
diffuse tenderness | 0
atrial fibrillation with rapid ventricular rate | 0
elevated white blood count | 0
ProBNP of 11,442 pg/mL | 0
negative COVID-19 test | 0
creatinine of 1.84 mg/dL | 0
elevated D-dimer of 6.45 mg/L | 0
minimal infiltrates | 0
cardiomegaly | 0
mild pleural effusion bilaterally | 0
normal ejection fraction | 0
no right heart strain | 0
right lower lobe pulmonary embolism | 0
mild abdominal ascites | 0
antibiotic coverage | 0
admitted to the intensive care unit | 0
urine and blood cultures drawn | 0
no micro-organisms | 0
abdominal discomfort | 24
afib RVR managed | 24
anticoagulated for PE | 24
paracentesis | 24
abdominal ultrasound-guided paracentesis | 24
4250 cc of dark straw-colored fluid | 24
ascitic fluid analysis | 24
no evidence suggestive of spontaneous bacterial peritonitis | 24
preliminary ascitic fluid pathology | 24
atypical epithelioid cells | 24
reactive mesothelial cells | 24
viral hepatitis serologies | 24
liver function tests | 24
Alpha-fetoprotein | 24
CA 19-9 | 24
CEA | 24
ANA | 24
anti-smooth muscle antibody | 24
anti-mitochondrial antibody | 24
noncontributory | 24
serum ascites albumin gradient | 24
SAAG of 0.8 | 24
new-onset nausea | 168
new-onset vomiting | 168
new-onset diarrhea | 168
repeat CT abdomen/pelvis | 168
multiple dilated loops of the small bowel | 168
high-grade small bowel obstruction | 168
thickened omentum | 168
questionable peritoneal carcinomatosis | 168
expedited to the operating room | 168
exploratory laparotomy | 168
extensive spread of the disease | 168
biopsies collected | 168
advanced carcinomatosis | 168
matted visceral structures | 168
probable malignant ascites | 168
rapidly decompensated | 360
expired | 360
final pathology report | 360
primary MPM | 360
abdominal fluid | 360
scattered and markedly atypical mesothelial cells | 360
suspicious for malignant mesothelioma | 360
mixed inflammation | 360
numerous histiocytes | 360
immunohistochemistry | 360
mesothelial phenotypic expression | 360
peritoneum excision | 360
malignant epithelioid mesothelioma | 360
rhabdoid features | 360