38 years old | 0\
male | 0\
HBV-associated PAN | -6 months\
acute abdomen | 0\
septic shock | 0\
prednisolone | -6 months\
cyclophosphamide | -6 months\
Tenofovir | -6 months to -2 months\
chronic renal failure | -6 months\
diabetes mellitus Type II | -6 months\
free sub diaphragmatic air | 0\
peritonitis | 0\
perforations of the small intestine | 0\
segmental enterectomy with anastomosis | 0\
mechanical ventilation | 0\
circulatory support | 0\
acute-on-chronic renal failure | 0\
weaned off the ventilator | 72\
haemodynamically stable | 72\
tenofovir | 72\
IV methylprednisolone | 72\
abdominal drain catheter presented enteric content | 168\
second explorative laparotomy | 168\
new perforations | 168\
multiple areas of patchy necrosis | 168\
suture repaired | 168\
open abdomen | 168\
plasma exchanges | 168\
IV cyclophosphamide | 168\
IV methylprednisolone | 168\
IV prednisone | 168\
third laparotomy | 240\
new necrotic lesions | 240\
suture repaired | 240\
necrotic lesion on the left lobe of the liver | 240\
fourth laparotomy | 336\
segmental enterectomy with anastomosis | 336\
cholecystectomy | 336\
anastomotic leak | 336\
gangrenous gallbladder | 336\
died | 360\
weight loss | -12 months\
myalgias | -12 months\
fever | -12 months\
skin erythema | -12 months\
deterioration of renal function | -12 months\
new onset of diabetes mellitus Type II | -12 months\
hypertension | -12 months\
HBsAg | 0\
HBeAg | 0\
Anti-HBcAb | 0\
absence of Anti-HBsAb | 0\
absence of Anti-HBeAb | 0