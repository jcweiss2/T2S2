63 years old | 0
woman | 0
two-day history of general body malaise | 0
two-day history of diarrhea | 0
two-day history of vomiting | 0
two-day history of influenza-like symptoms | 0
admitted to the hospital | 0
increased confusion | 0
splenectomy 43 years earlier | -376968
idiopathic thrombocytopenic purpura | -376968
menometrorrhagia | -376968
vaccinated with PPV23 | -376968
antibody response tested | -672
antibody response adequate | -672
fever | 0
hypotension | 0
bradycardia | 0
tachypnea | 0
decreased oxygen saturation | 0
cyanosis of the lips | 0
cyanosis of the distal extremities | 0
no neck stiffness | 0
no meningeal reactions | 0
normal cardiac auscultation | 0
normal pulmonic auscultation | 0
soft abdomen | 0
non-tender abdomen | 0
diagnosed with severe sepsis | 0
volume therapy started | 0
blood cultures | 0
broad-spectrum antimicrobial therapy started | 0
cefuroxim | 0
gentamicin | 0
metronidazole | 0
hydrocortisone | 0
white blood cell count elevated | 0
neutrophils elevated | 0
hemoglobin low | 0
thrombocytes low | 0
CRP elevated | 0
P-lactate elevated | 0
aB-P-O2 elevated | 0
aB-P-CO2 low | 0
aB-pH elevated | 0
Streptococcus pneumococcal urinary antigen positive | 0
chest x-ray pulmonic stasis | 0
transferred to ICU | 24
disseminated intravascular coagulation | 24
microthrombi in hands | 24
microthrombi in feet | 24
blood cultures grew S. pneumoniae | 48
antimicrobial therapy changed to penicillin G | 48
MIC <0.1 μg/ml | 48
suspicion of endocarditis | 72
TTE performed | 72
TTE showed hypokinesia | 72
ejection fraction 45% | 72
endocarditis dismissed | 72
necrosis of fingertips | 72
necrosis of toes | 72
renal insufficiency | 72
hemodialysis started | 72
antibiotic therapy changed to ceftriaxone | 72
leucocytes decreased | 96
CRP decreased | 96
fever resolved | 96
tracheal secret culture negative | 96
transferred to medical department | 216
antibiotics stopped | 216
serotype 12F identified | 216
afebrile | 264
fluctuating CRP | 264
condition improved | 264
discharged | 528
oral dicloxacillin prescribed | 528
raised leucocytes | 528
raised CRP | 528
suspected infection site necrotic tissue | 528
wound cultures S. aureus | 528
wound cultures haemolytic streptococci group C/G | 528
TTE unchanged | 528
necrotic fingers amputated | 2232
necrotic toes amputated | 2232
readmitted with severe sepsis | 3720
sepsis regimen started | 3720
ceftriaxone therapy started | 3720
TEE performed | 3720
endocarditis diagnosed | 3720
moving elements on aortic valve | 3720
blood cultures grew S. pneumoniae | 3720
antimicrobial therapy changed to penicillin G | 3720
MIC <0.1 μg/ml | 3720
treated conservatively with penicillin G | 3720
recovered | 3720
serotype 12F identified | 3720
serological tests performed | -15672
antibody levels sufficient | -15672
antibody levels tested 18 months before first IPD | -15672
antibody levels tested between IPD episodes | 2640
antibody levels tested 1 year after second IPD | 8760
antibodies to 12F present | -15672
antibodies to 12F present | 2640
antibodies to 12F present | 8760
