47 years old | 0
female | 0
admitted to the hospital | 0
postoperative bleeding | -24
vaginal hysterectomy | -24
third-degree uterovaginal prolapse | -24
conscious but drowsy | 0
tachypneic | 0
heart rate 120 beats per minute | 0
blood pressure 90/60 mm Hg | 0
peripheries cold and clammy | 0
low hemoglobin 6.2 g/dl | 0
emergency laparotomy | 0
triple lumen central venous access | 0
fluid resuscitation | 0
inotropic support | 0
left radial artery cannulation | 0
invasive hemodynamic monitoring | 0
surgery | 0
ligation of bilateral internal iliac arteries | 0
intraoperative fresh frozen plasma | 0
intraoperative packed red blood cells | 0
inotropic support with dopamine | 0
admitted in intensive care unit | 0
elective ventilation | 0
disseminated intravascular coagulopathy | 48
blood products | 48
cryoprecipitate | 48
inotropic support with dopamine | 48
acute respiratory distress syndrome | 72
increasing ventilatory support | 72
tracheostomy | 168
ventilatory support | 168
dusky discoloration of the digits | 72
cold extremities | 72
deferred decannulation | 72
worsening of discoloration | 120
left radial artery cannula removal | 120
vascular surgery opinion | 120
Doppler ultrasound | 120
partial thrombosis | 120
injection Clexane | 120
IV low molecular weight Dextran | 120
stellate ganglion block | 120
nitroglycerine ointment | 72
discoloration improvement in right hand | 120
discoloration worsening in left hand | 120
dry gangrene | 192
pulmonary rehabilitation | 720
psychiatric rehabilitation | 720
amputation of gangrenous digits | 720
brachial plexus block | 720