33 years old | 0
man | 0
admitted to the hospital | 0
severe anemia | 0
unresponsive to hemotransfusions | 0
increasing doses of erythropoietin | 0
membranoproliferative glomerulonephritis | -43824
renal biopsy | -43824
steroids | -43824
immunosuppressants | -43824
persistent proteinuria | -43824
microhematuria | -43824
glomerular sclerosis | -43824
mesangiocapillary global proliferation | -43824
fibrinoid necrosis | -43824
vascular thrombosis | -43824
extracapillary proliferation | -43824
Congo red staining for amyloid | -43824
immunofluorescence (IF) results | -43824
tiny granular deposits | -43824
semilinear membrane for immunoglobulin G (IgG) | -43824
C3 | -43824
immunoglobulin A (IgA) | -43824
immunoglobulin M (IgM) | -43824
C1q | -43824
κ and λ light chains | -43824
accumulation of intravascular fibrinogen | -43824
azathioprine | -43824
mycophenolate | -43824
steroid therapy | -43824
rapid reduction in proteinuria | -43824
disappearance of microhematuria | -43824
bilateral aseptic necrosis of the femoral head | -26208
stopped steroids | -17520
slow worsening renal function | -17520
serum creatinine: 2.5 mg/dL | -17520
proteinuria (1.5-2 g/24 h) | -17520
anemia | -17520
darbepoetin alfa | -17520
admitted to the emergency room | -72
hospitalized | 0
severe anemia (hemoglobin: 6 g/dL) | 0
severe asthenia | 0
dyspnea even for minor efforts | 0
hemoglobin values increased after hemotransfusion | 0
colonoscopy | 0
gastroscopy | 0
peripheral smear | 0
schistocytes | 0
direct Coombs tested negative | 0
indirect Coombs tested negative | 0
G6PDH appeared within the normal range | 0
haptoglobin reduced | 0
lactate dehydrogenase increased slightly | 0
direct bilirubin levels normal | 0
indirect bilirubin levels normal | 0
autoimmunity normal | 0
persistent slight reduction in C3 | -52560
hemoglobin levels decreased by 7 g/dL | 72
infusion of a new unit of packed red blood cells | 72
full-abdomen ultrasound scan | 72
blood abdominal collections | 72
significant changes | 72
kidney size reduction | 72
chest X-ray imaging | 72
bronchopneumonia bilaterally spread in the middle lobe | 72
hemoptysis with bright red blood and clots | 96
coughing for several days | 96
chest computed tomographic (CT) scan | 96
multilobar alterations extended to both lungs | 96
ground-glass appearance | 96
intralobular involvement | 96
intra-acinar involvement | 96
thickening of the interlobular septa | 96
distortion and rails and interlobular fissures | 96
Diffusion lung CO (DLCO) analysis | 96
increase in DLCO (157%) | 96
reduction in alveolar volume | 96
intra-alveolar hemorrhage | 96
methylprednisolone | 96
prednisone 1 mg/kg/d | 96
azathioprine | 96
low-flow oxygen therapy | 96
anti-glomerular basement membrane (anti-GBM) antibodies | 96
false-negative serum cases | 96
IF | 96
chemiluminescence | 96
C-ANCA | 96
P"|ANCA | 96
transnasal endoscopy | 96
bleeding striae in the first tracheal rings | 96
bronchoscopy | 120
lesions visible at tracheal level | 120
bronchoalveolar lavage was blood | 120
fibrinoid necrosis | 120
improvement in the clinical picture | 144
test results | 144
fatigue | 144
dyspnea gradually reduced | 144
oxygen saturation progressed satisfactorily | 144
further transfusions | 144
peripheral oxygen saturation maintained at around 98% | 144
deterioration of renal function | 168
filtrate of 17 mL/min reduced to 11 mL/min | 168
increase in blood urea | 168
increase in creatinine values | 168
increase in potassium concentrations | 168
increase in phosphorus concentrations | 168
peritoneal dialysis | 168
CT control chest | 480
improvement in both lungs | 480
thickening of the bronchial walls | 480
interlobular septa persisted | 480
spirometry | 480
DLCO test | 480
immunosuppressive therapy reduced | 480
discharged | 480
hemoglobin level maintained | 480
erythropoiesis-stimulating agent doses | 480
automated peritoneal dialysis | 480
suspension of immunosuppressive therapy | 1296
dosage of Ab anti-GBM | 1296
negative antibodies | 1296
