66 years old | 0
male | 0
admitted to the hospital | 0
COVID-19 infection | 0
hypertension | -25920
angiotensin-converting-enzyme inhibitor | -25920
diabetes | -62496
metformin 850 mg/d | -62496
HbA1c 6.3% | -62496
acute respiratory failure | 0
hemodynamically stable | 0
neurologically stable | 0
dyspneic | 0
respiratory rate 25/min | 0
oxygen saturation SpO2% 83% | 0
temperature 39.7°C | 0
weight 99 kg | 0
height 1.76cm | 0
body mass index 31.96kg/m2 | 0
unremarkable clinical examination | 0
RT-PCR for SARS-COV 19 positive | 0
nonenhanced chest CT scan showing peripheral ground-glass opacities | 0
pulmonary involvement 25% to 50% | 0
lymphopenia | 0
increased ferritin | 0
increased CRP | 0
increased LDH | 0
hypoxemia | 0
Partial Pressure of Oxygen 55 mm Hg | 0
hospitalized in intensive care unit | 0
oxygen therapy via nasal cannula 7l/min | 0
SpO2% 93% | 0
difficulty in breathing | 72
SpO2 decreased to 84% | 72
severe hypoxemia | 72
Partial Pressure of Oxygen 47 mm Hg | 72
contrast-enhanced chest CT showing worsening pulmonary involvement | 72
pulmonary involvement more than 75% | 72
oxygen therapy with high-concentration mask 14l/min | 72
prone decubitus sessions | 72
SpO2 90% | 72
favorable evolution | 72
sudden onset of palpitations | 120
worsening dyspnea | 120
heart rate 186 bpm | 120
blood pressure 134/80 mm Hg | 120
atrial fibrillation | 120
rhythm control strategy | 120
amiodarone continuous infusion | 120
amiodarone initial bolus | 120
HR slowed | 120
HR not dropping below 140 bpm | 120
new atrial fibrillation | 122
ventricular response 205 bpm | 122
hemodynamic instability | 122
BP 70/50 mm Hg | 122
altered state of consciousness | 122
Glasgow Coma Scale 8/15 | 122
external electric shock 260J | 122
sinus rhythm restored | 122
HR 98 bpm | 122
hemodynamically stabilized | 122
BP 125/80 mm Hg | 122
no recovery of normal consciousness | 122
suspected stroke | 122
cerebral MRI | 123
brainstem acute ischemic stroke | 123
National Institutes of Health Stroke Scale score 35 | 123
contraindicated thrombolysis | 123
severe neuro0vegetative disorders | 123
prolonged apnea | 123
extreme bradycardia | 123
tachycardia | 123
unrecovered cardiac arrest | 125
refractory ventricular fibrillation | 125
resuscitation measures | 125
