32 years old | 0
female | 0
admitted to the ICU | 0
severe coronavirus disease 2019 | 0
hypoxemic respiratory failure | 0
SpO2: 94% with oxygen therapy | 0
respiratory rate of 30 breaths per min | 0
piperacillin–tazobactam | 0
methylprednisolone | 0
remdesivir | 0
high-flow nasal cannula therapy | 0
intubated | 0
standard lung-protective ventilation | 0
pregnancy terminated | 0
acute respiratory distress syndrome worsening | 0
nonstress test revealed fetal distress | 0
lower segment cesarean section | 0
live female baby delivered | 0
PaO2/FiO2 ratio post LSCS was 120 | 0
two prone ventilation sessions | 0
significant improvement in oxygenation | 0
P/F Ratio to 300 | 0
diffuse subcutaneous edema of the face | 0
subcutaneous edema reduced over next 4 days | 96
percutaneous tracheostomy | 168
septic shock with Klebsiella pneumoniae bacteremia | 168
antimicrobials as per sensitivity report | 168
colistin | 168
meropenem | 168
shock recovered | 168
weaning initiated | 384
spontaneous breathing trial | 384
inability to close left eyelid | 384
deviation of angle of mouth to the right side | 384
no other focal neurological deficit | 384
plantar reflexes flexor response | 384
examination of ears showed no discharge | 384
power of all four limbs reduced | 384
Medical Research Council sum score of 40 | 384
critical illness neuromyopathy | 384
patching of eyelid | 384
lubrication with eye drops | 384
contrast-enhanced computed tomography scan | 384
soft-tissue swelling with fat stranding in left cheek and masseter muscle | 384
no evidence of stroke | 384
no significant compression in tract of facial nerve | 384
no fracture or osseous lesion in facial canal | 384
active limb physiotherapy | 384
good glycemic control | 384
steroids deferred | 384
acyclovir not administered | 384
weaned from mechanical ventilation | 552
decannulated | 720
left facial nerve palsy persisted | 720
House–Brackmann Facial Nerve Grade IV | 720
magnetic resonance imaging of the brain | 720
subtle postcontrast enhancement in cisternal and intracanalicular part of 7th and 8th nerve complex | 720
discharged home | 720
eye care instructions | 720
complete resolution of paresis | 2160
no long-term effects | 2160
