23 years old | 0
    woman | 0
    presented with sore throat | 0
    nausea | 0
    subjective fever | 0
    chills | 0
    sore throat | -24
    oral antibiotics | -24
    febrile | 0
    temperature of 102.2° Fahrenheit | 0
    tachycardic | 0
    heart rate of 130 beats per minute | 0
    hypotensive | 0
    blood pressure of 90/50 mm Hg | 0
    leukocyte count of 17.87 k/ul | 0
    predominant neutrophil count of 86.8% | 0
    elevated creatinine of 3.6 mg/dL | 0
    sepsis | 0
    acute kidney injury | 0
    empiric antibiotics | 0
    rapid crystalloid infusion | 0
    hypotensive persisted | 0
    admitted to intensive care unit | 0
    fulminant septic shock | 0
    Streptococcus anginosus isolated from blood cultures | 0
    Fusobacterium necrophorum isolated from blood cultures | 0
    computed tomography of the chest | 0
    scattered bilateral nodular opacities | 0
    peripheral distribution suspicious for septic emboli | 0
    small bilateral pleural effusions | 0
    adjacent consolidations | 0
    empiric piperacillin/tazobactam | 0
    metronidazole | 0
    Lemierre's syndrome suspected | 0
    internal jugular vein thrombosis ruled out | 0
    computed tomography of the neck | 0
    repeat computed tomography of the chest | 240
    decrease in size of bilateral nodular opacities | 240
    new areas of cavitation | 240
    increased moderate left pleural effusion | 240
    near complete atelectasis of left lower lobe | 240
    left sided chest tube placed | 240
    parapneumonic effusion | 240
    F. necrophorum sensitive to augmentin | 0
    F. necrophorum sensitive to clindamycin | 0
    F. necrophorum sensitive to imipenem | 0
    F. necrophorum resistant to metronidazole | 0
    Streptococcus anginosus pansensitive to penicillin | 0
    Streptococcus anginosus pansensitive to ceftriaxone | 0
    Streptococcus anginosus pansensitive to clindamycin | 0
    Streptococcus anginosus pansensitive to vancomycin | 0
    Streptococcus anginosus pansensitive to levofloxacin | 0
    Streptococcus anginosus pansensitive to erythromycin | 0
    antibiotics switched to piperacillin/tazobactam | 0
    antibiotics switched to clindamycin | 0
    diagnosed with Lemierre's syndrome | 0
    secondary to F. necrophorum | 0
    pulmonary septic emboli | 0
    stay of 18 days in hospital | 432
    clinical condition improved | 432
    discharged home | 432
    ceftriaxone | 432
    clindamycin | 432
    outpatient follow-up | 432
    good recovery | 432
