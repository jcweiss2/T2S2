71 years old | 0
female | 0
admitted to the emergency department | 0
complaint of a painful abdominal mass | 0
malnourished | 0
poor hygiene | 0
febrile | 0
temperature of 38℃ | 0
pulse rate was 106 beats per minute | 0
no evidence of a heart murmur | 0
no lung crackles on auscultation | 0
breath sounds were clear | 0
no signs of abdominal or rebound tenderness | 0
large tender mass in the abdominal left upper quadrant | 0
hemoglobin, 8.3 g/dl | 0
white blood cell count, 17,510/ml | 0
blood urea nitrogen, 27.5 mg/dl | 0
creatinine, 0.38 mg/dl | 0
sodium, 142 mEq/L | 0
chloride, 105 mEq/L | 0
potassium, 3.2 mEq/L | 0
C-reactive protein, 304 mg/L | 0
urinalysis revealed no abnormalities | 0
chest radiography showed no abnormalities | 0
computed tomography of the abdomen revealed a large abscess pocket | 0
incised the mass and drained a large abscess | 0
diagnostic laparotomy | 0
gastric cancer invading the abdominal wall | 0
no apparent distant metastasis | 0
peritoneal cavity was not contaminated | 0
dissection of the stomach from the peritoneal membrane was impossible | 0
total gastrectomy along with resection of the involved abdominal wall | 0
resection of peritoneum, rectus abdominis muscle, and subcutaneous tissue | 0
no remaining muscle or subcutaneous layer on the patient's left upper quadrant | 0
overlying skin was not viable | 0
wet gauze packing of the wound | 0
D1 lymph node dissection for the perigastric lymph nodes | 0
hypotensive | 0
septic | 0
R status was expected to be R1 | 0
admitted to the intensive care unit | 0
postoperative care | 0
resuscitation | 0
vital signs became stable on the first postoperative day | 24
febrile with a temperature of 38.8℃ on the first postoperative day | 24
chest radiography showed diffuse haziness in both lung fields on the first postoperative day | 24
suspicion of pneumonia | 24
intensive treatment, including broad-spectrum antibiotics and parenteral nutrition | 24
closely observed for suspicious leakage at the anastomosis | 24
resumed oral intake on the third postoperative day | 72
chest radiography on the seventh postoperative day showed improvement of the pneumonia | 168
moved to a general ward on the eighth postoperative day | 192
resumed ambulation on the eighth postoperative day | 192
wet dressing of the wound | 192
abdominal binder was used to prevent evisceration | 192
planned to perform chemotherapy | 192
growth of the cancer progressed rapidly | 960
wound had filled with growing cancer on the 40th postoperative day | 960
prognosis was expected to deteriorate | 960
conservative management, including analgesics, sedatives, and nutrition for palliation | 960
oral intake was impossible on the 60th postoperative day | 1440
intestinal obstruction on the 60th postoperative day | 1440
died of multiorgan failure caused by sepsis and pneumonia on the 82nd postoperative day | 1968
histologic diagnosis was poorly differentiated adenocarcinoma of the stomach | 1968
13 lymph nodes harvested, 5 were cancer-cell positive | 1968
N2 | 1968
T stage could not be determined | 1968
suspected to be T4a | 1968
cancer stage was IIIB | 1968