62 years old | 0
female | 0
presented with necrotizing fasciitis of left thigh and groin | 0
carbuncle | -336
chills | -336
no pyrexia | -336
diet-controlled type 2 diabetes mellitus | 0
hemoglobin A1c level 5.7% | 0
ascorbic acid 1,000 mg daily | 0
denied non-steroidal anti-inflammatory drugs | 0
denied smoking | 0
denied illicit drug use | 0
alcohol consumption | 0
hypotensive | 0
blood pressure 87/63 mm Hg | 0
pulse 92 bpm | 0
temperature 36.6°C | 0
severe tenderness left thigh | 0
posterior crepitus | 0
intravenous fluid resuscitation | 0
urgent imaging | 0
hemoglobin 7.8 g/dl | 0
mean corpuscular volume 71.9 fl | 0
white blood cell count 11.9 × 103 µl | 0
platelet count 151 × 103 µl | 0
reticulocyte count 3.39% | 0
immature reticulocyte fraction 35.80% | 0
serum iron level 7.0 µg/dl | 0
serum transferrin level 123 mg/dl | 0
total iron-binding capacity 7.0 µg/dl | 0
negative Direct Coombs test | 0
negative fecal occult blood testing | 0
CT scan showing air in posterior thigh muscles | 0
air extending to gluteus maximus | 0
air extending to knee | 0
indicative of necrotizing fasciitis | 0
started on intravenous vancomycin | 0
started on clindamycin | 0
started on piperacillin/tazobactam | 0
aggressive fluid resuscitation for septic shock | 0
fasciotomy | 0
debridement | 0
extensive devitalized tissue | 0
necrosis left thigh | 0
disarticulation left lower extremity | 0
intraoperative wound culture grew C. septicum | 0
managed in intensive care unit | 0
screening colonoscopy planned in 2 months | 0
antibiotic regimen changed to clindamycin | 0
antibiotic regimen changed to piperacillin/tazobactam | 0
frank blood in fecal management tube | 288
emergent colonoscopy | 288
fungating polypoid mass in cecum | 288
sessile mass | 288
ulcerated mass | 288
partially obstructing mass | 288
histopathology consistent with invasive adenocarcinoma | 288
laparoscopic right hemicolectomy | 432
CT imaging negative for metastatic spread | 432
no signs or symptoms of recurrence of colon cancer | 0
Clostridium septicum infection | 0
association with colon cancer | 0
negative metastatic spread | 0
limb amputation | 0
discharge after treatment | 0
outpatient follow-up | 0
