62 years old | 0
male | 0
non-smoker | 0
presented to the emergency department | 0
worsening pain in the left groin | -672
subjective fevers | -672
ChAdOx1 nCoV-19 vaccine second dose | -336
episode of diarrhoea | -240
no recent history of taking antibiotics | 0
total replacement of the left hip | -131400
arthrosis secondary to hip dysplasia | -131400
minor asymptomatic osteolysis secondary to metal-on-metal wear | -131400
hypertension | 0
paroxysmal atrial fibrillation | 0
rivaroxaban | 0
admitted to a hospital six years prior | -52560
diarrhoea | -52560
haematochezia | -52560
Bacteroides vulgatus bacteremia | -52560
inpatient gastroscopy | -52560
colonoscopy | -52560
full recovery | -52560
no significant gastrointestinal abnormality | -52560
no risk factors for immunocompromise | 0
afebrile | 0
mild tachycardia | 0
heart rate of 100-110 bpm in atrial fibrillation | 0
hypotensive | 0
blood pressure of 80/40 mmHg | 0
respiratory rate of 19 breaths per minute | 0
SpO2 99% on room air | 0
left hip joint irritability to passive movements | 0
cardiovascular findings unremarkable | 0
gastrointestinal findings unremarkable | 0
respiratory findings unremarkable | 0
elevated levels of inflammatory markers | 0
normal blood metal ion levels | 0
pelvic x-ray showed no new changes to the prosthesis | 0
longstanding femoral osteolysis secondary to metal wear | 0
aspiration of the hip yielded 20 mL haemoserous fluid | 0
white blood cell count 250,200 WBC/µL | 0
gram-negative bacilli detected | 0
gram-positive bacilli detected | 0
started on empirical intravenous cefazolin | 0
transferred to intensive care unit | 0
light growth of tiny, grey, translucent colonies on day 2 | 48
identified as F. plautii on day 4 | 96
MALDI-TOF MS confirmation | 96
growth in peripheral blood culture anaerobic bottle | 96
antibiotic regimen changed to amoxycillin-clavulanate, gentamicin, metronidazole, vancomycin | 96
antibiotic susceptibility determined on day 4 | 96
surgical intervention delayed due to COVID-19 | 96
medical stabilisation in intensive care unit | 96
first-stage revision hip arthroplasty on day 7 | 168
exploration of hip via posterior approach | 168
extensive abscess formation | 168
destruction of soft tissue deep to the fascia | 168
no gross evidence of metalosis | 168
no loosening of the stem | 168
use of fine oscillating saw | 168
good fixation of acetabular component | 168
use of Explant® acetabular cup removal system | 168
debridement of pericapsular soft tissue erosion | 168
pulse lavage | 168
intermittent irrigation with hydrogen peroxide | 168
reaming of the canal with 14 mm flexible reamer | 168
thorough washing with canal brush | 168
extraction of all hardware | 168
implantation of antibiotic cement articulating spacer | 168
no organisms isolated on intraoperative culture | 168
thickened ascending colon on CT abdomen | 168
colonoscopic biopsy showed sigmoid tubular polyp | 168
diverticular disease | 168
conservative management | 168
normal chest x-ray | 168
normal uranalysis | 168
normal cardiac echocardiogram | 168
ceftriaxone 2 g intravenously for six weeks | 168
oral amoxicillin/clavulanic acid and metronidazole for six weeks | 168
normalisation of C-reactive protein | 168
further aspiration of the hip | 168
yielded 832 WBC/µL | 168
20% polymorphonuclear cells | 168
negative cultures | 168
second stage revision arthroplasty three months after first stage | 2160
posterior approach for exposure | 2160
extraction of antibiotic cement | 2160
extraction of spacer implants | 2160
no macroscopic evidence of infection | 2160
no bone necrosis | 2160
multiple swabs and tissue cultures negative | 2160
administration of intraoperative cefazolin and vancomycin | 2160
preparation of acetabular and femoral sides | 2160
implantation of uncemented components | 2160
discharged on day 7 | 2160
uncomplicated recovery | 2160
at 12-month follow-up in good health | 2160
no ongoing infective issues | 2160
off antibiotics | 2160
normal, pain-free gait | 2160
near normal hip range of movement | 2160
