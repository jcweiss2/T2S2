65 years old|0
female|0
presented with right flank pain|-168
presented with fatigue|-168
immobile at home|-24
transported by ambulance|-24
diabetes mellitus|0
breast cancer|-87600
Glasgow Coma Scale: E4V5M6|0
blood pressure 77/55 mm Hg|0
heart rate 120 beats/min|0
temperature 36.2°C|0
respiratory rate 42/min|0
mildly distended abdomen|0
right flank tenderness|0
costovertebral angle tenderness|0
white blood cell count 18.5x10^9/L|0
hemoglobin 11.7 × 10^-1 g/L|0
platelet 7.8×10^-5/L|0
blood urea nitrogen 67.9 mg/dL|0
creatinine 3.53 mg/dL|0
sodium 124 mEq/L|0
potassium 3.7 mEq/L|0
chloride 84 mEq/L|0
prothrombin time-international normalized ratio 1.29|0
blood glucose 543 mg/dL|0
glycosylated hemoglobin A1c 12.1%|0
metabolic acidosis|0
pH 7.41|0
arterial oxygen pressure 101.6 mm Hg|0
PaCO2 16.1 mm Hg|0
bicarbonate 10.0 mEq/L|0
base excess 12.1 mEq/L|0
lactic acid 3.43 mmol/dL|0
urinalysis white blood cell 3+|0
urinalysis occult blood 3+|0
CT scan emphysematous changes in right kidney|0
diagnosis of right emphysematous pyelonephritis class 3B|0
admitted to ICU|0
blood cultures obtained|0
urine cultures obtained|0
meropenem administered intravenously|0
vancomycin administered intravenously|0
resuscitation with intravenous fluids|0
resuscitation with vasopressors|0
resuscitation with steroids|0
condition deteriorated|0
intubated|6
mechanical ventilation required|6
portable abdominal X-ray progression of emphysematous changes|6
exploratory laparotomy|6
swelling in Gerota’s fascia|6
release of foul-smelling gas|6
spongy renal parenchyma|6
purulent material drained|6
right nephrectomy performed|6
copious irrigation|6
abdomen closed|6
returned to ICU postoperatively|6
cultures revealed Escherichia coli|6
antibiotics continued for 14 days|6
leukocytosis subsided|168
fever subsided|168
acute renal failure postoperatively|6
hemodialysis required|6
tracheostomy performed|6
prolonged mechanical ventilation required|6
weaned from hemodialysis|168
weaned from mechanical ventilation|168
transferred to rehabilitation hospital|504
