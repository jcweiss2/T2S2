66 years old | 0
male | 0
diabetes mellitus | -10080
benign prostatic hyperplasia | -10080
fatigue | -504
suprapubic tenderness | -72
urinalysis | -72
protein 1+ | -72
glucose 3+ | -72
blood 3+ | -72
no nitrites | -72
no leukocyte esterase | -72
ultrasound | -72
moderate hydronephrosis | -72
urinary retention | -72
Foley catheter | -72
2.3 L of urine | -72
improved symptoms | -72
lethargy | -168
hyperglycemia | -168
blood glucose 840 mg/dL | -168
dysuria | -168
urine culture positive for E. coli | -168
blood culture positive for E. coli | -168
hemoglobin A1c 13.6% | -168
computed tomography | -168
extensive gas within bilateral renal parenchyma | -168
gas within left renal sinus | -168
perinephric fat stranding | -168
thickening of Gerota's fascia | -168
septic shock | 0
bilateral radical nephrectomy | 0
dialysis-dependent | 24
readmitted | 168
recurrent MDR E. coli pyocystitis | 168
anemia | 168
persistent urinary retention | 168
intravenous antibiotics | 168
red blood cell transfusions | 168
iron supplementation | 168
suprapubic catheter placement | 168
emphysematous pyelonephritis | 0
bilateral emphysematous pyelonephritis | 0
multifocal hemorrhage | 0
acute pyelonephritis | 0
abscesses | 0
infarction | 0
gas-filled cysts | 0
vasculitis | 0
diabetic nephropathy | -10080
diffuse thickening of glomerular and tubular basement membranes | -10080
mesangial expansion | -10080
diffuse acute tubular injury | 0
loss of proximal tubule brush border | 0
simplified tubular epithelium | 0
sloughed epithelial cells | 0
mild-to-moderate intimal fibrosis | 0
arteriosclerosis | 0
thickening of arteriolar walls | 0