64 years old | 0
female | 0
bipolar depression | 0
diabetes | 0
migraine headaches | 0
seizure disorder | 0
admitted to the hospital | 0
found unresponsive | -1
ambient temperature over 90°F | -1
amitriptyline 175 mg daily | -672
cyclobenzaprine 10 mg daily | -672
lurasidone 80 mg daily | -672
benztropine 1 mg three times a day | -672
topiramate extended release 100 mg daily | -672
clonazepam 0.5 mg daily | -672
trazodone 100 mg daily | -672
sitagliptin 25 mg daily | -672
erenumb 70 mg injected monthly | -672
febrile | -1
emergency medical service called | -1
cool compresses applied | -1
transported to the hospital | -1
hypotensive | 0
blood pressure 84/42 | 0
rectal temperature 42°C | 0
skin warm and dry | 0
mucous membranes dry | 0
responsive to painful stimuli | 0
leucocytosis | 0
creatinine phosphokinase normal | 0
EKG normal | 0
admitted to ICU | 0
started on vancomycin | 0
started on cefepime | 0
blood cultures grew Staphylococcus hominis | 24
core body temperature decreased | 24
mentation returned to baseline | 24
transferred to medical floor | 48
treated for Staph hominis bacteraemia | 48
7-day course of vancomycin | 48
discontinued cyclobenzaprine | 120
feeling overheated and fatigued for 2 weeks | -336
follow-up call | 1440
primary care physician advised to continue medication regimen | 1440
educated about risks of polypharmacy | 1440
discussed medication changes | 1440