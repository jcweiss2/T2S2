84 years old | 0
male | 0
admitted to the hospital | 0
lethargy | -72
fatigue | -72
weakness | -72
bloody urine | -24
intermittent fevers | -24
ischemic cardiomyopathy | 0
heart failure | 0
atrial fibrillation | 0
taking Coumadin | 0
lived in Upstate New York | 0
hepatosplenomegaly | 0
petechial rash | 0
elevated total bilirubin | 0
elevated alkaline phosphatase | 0
elevated AST | 0
elevated ALT | 0
elevated INR | 0
low albumin | 0
low hemoglobin | 0
low platelet count | 0
ascites | 0
CBD diameter of 0.5 cm | 0
given fresh frozen plasma | 24
given vitamin K | 24
intermittent fevers | 24
blood cultures negative | 24
increasing bilirubin | 24
paracentesis | 120
low ascites albumin | 120
low serum albumin | 120
high neutrophil count in ascites fluid | 120
low haptoglobin | 120
worsening encephalopathy | 120
hypotensive | 120
transferred to ICU | 120
peripheral smear obtained | 120
intraerythrocytic organisms seen | 120
initiation of intravenous clindamycin | 120
initiation of quinine | 120
increasing bilirubin | 144
serum serology for Lyme negative | 144
serum serology for Erlichia negative | 144
serum serology for anaplasmosis negative | 144
patient passed away | 168