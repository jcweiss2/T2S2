25-year-old | 0  
    primigravida | 0  
    pregnancy | 0  
    uncomplicated | 0  
    well before delivery | 0  
    hospital attendance | 0  
    spontaneous onset of labor | 0  
    fetal distress | -2  
    second stage of labor | -2  
    ventouse-assisted delivery | -1  
    male infant born | 0  
    birth weight 3940 grams | 0  
    immediate resuscitation | 0  
    mask ventilation | 0  
    intubated | 8  
    poor respiratory effort | 8  
    transferred to NICU | 8  
    SIPPV | 8  
    minimal pressures | 8  
    no additional oxygen requirement | 8  
    empirical antibiotics | 8  
    early-onset sepsis | 8  
    gentamicin | 8  
    benzyl penicillin | 8  
    respiratory support weaned | 13.5  
    extubated | 13.5  
    neutropenia | 18  
    left shift | 18  
    CRP elevated | 18  
    procalcitonin elevated | 18  
    lumbar puncture | 23  
    normal cell count | 23  
    negative for pathogens | 23  
    placental eSwab | 23  
    pure growth | 23  
    Gram-negative diplococci | 23  
    MALDI-TOF | 23  
    Neisseria meningitidis | 23  
    PCR ctrA | 23  
    PCR porA | 23  
    PCR serogroups | 23  
    serogroup W CC11 | 23  
    blood cultures negative | 29  
    heel-prick blood | 5.5  
    N. meningitidis DNA | 5.5  
    no maternal antibiotics | 0  
    funisitis | 23  
    chorioamnionitis | 23  
    ascending infection | 23  
    maternal inflammatory response | 23  
    fetal inflammatory response | 23  
    benzylpenicillin dosage decreased | 13.5  
    cefotaxime | 13.5  
    5-day course | 13.5  
    clinical improvement | 13.5  
    maternal leucocytosis | -2.5  
    neutrophil count elevated | -2.5  
    mother well postpartum | 0  
    baby discharged | 192  
    contact tracing | 192  
    chemoprophylaxis | 192  
    vaccination | 192  
    counseling | 192  

    