3 years old|0
female|0
dry cough|-336
gradual onset of dyspnea|-336
no fever|-336
no evidence of upper respiratory tract infection|-336
significant weight loss|0
progressive fatigue|0
chest X-ray showed heterogeneous opacity|0
pneumonia diagnosis|0
antibiotics (amoxicillin)|0
bronchodilators|0
cough not improved|0
dyspnea not improved|0
weakness of both lower limbs|-168
complete inability to walk|-168
flaccid weakness of lower limbs|-168
dyspnea persisted|0
admitted to local hospital|0
Guillain-Barré syndrome as differential diagnosis|0
condition worsened|0
dyspnea worsened|0
central cyanosis|0
referred to tertiary center|0
mechanical ventilation|0
severely dyspneic|0
respiratory rate 50 cycles/minute|0
SpO2 85%|0
loss of sphincter control|0
bladder palpable below umbilicus|0
catheterization|0
right-side supraclavicular lymph nodes|0
poor air entry in right lung|0
flaccid paraparesis|0
loss of tone|0
loss of reflexes|0
equivocal Babinski reflex|0
sensory examination inconclusive|0
opsoclonus-myoclonus eye movements|0
normal pupils|0
admitted to respiratory care unit|0
synchronized mechanical ventilation|0
serum electrolytes normal|0
unremarkable blood tests|0
respiratory acidosis|0
emergency chest MRI|0
large posterior-superior mediastinal mass|0
trachea deviation|0
pleural effusion|0
supraclavicular lymph nodes|0
dorsal spine invasion|0
canal stenosis|0
liver normal|0
whole-spine MRI|0
tumor extension to intraspinal canal|0
neuroblastoma differential diagnosis|0
high urine VMA|0
bone marrow biopsy confirmed neuroblastoma|0
thoracotomy|0
total resection of mass|0
spinal decompression|0
canal stenosis relief|0
pedicle screw instrumentation|0
histopathology: poorly differentiated neuroblastoma|0
supraclavicular lymph node biopsy|0
Shimada grading system|0
INRSS high-risk|0
postoperative improvement of dyspnea|0
weaning from ventilator|0
residual lower limb weakness|0
opsoclonus myoclonus eye movement|0
loss of bladder control|0
induction chemotherapy|0
cyclophosphamide|0
etoposide|0
vincristine|0
death due to pancytopenia|0
septicemia|0
renal impairment|0
intensive care|0
management|0
