59 years old | 0
male | 0
chronic obstructive pulmonary disease | 0
presented to the emergency department | 0
generalized fatigue | -72
dyspnea | -72
oliguria | -72
blood pressure 70/40 mmHg | 0
pulse rate 122 bpm | 0
temperature 36.4°C | 0
peripheral oxygen saturation 88% | 0
decreased breath sounds in lower right lung fields | 0
pretibial edema (++) | 0
hepatomegaly | 0
serum potassium 6.0 mEq/dL | 0
phosphorus 5.2 mg/dL | 0
alanine aminotransferase 672 U/L | 0
alkaline phosphatase 489 U/L | 0
total bilirubin 1.6 mg/dL | 0
direct bilirubin 0.87 mg/dL | 0
lactate dehydrogenase 2954 U/L | 0
creatinine 2.15 mg/dL | 0
uric acid 20.32 mg/dL | 0
serum calcium level 10.2 mg/dL | 0
albumin 3.0 g/dL | 0
C-reactive protein 115 mg/L | 0
chest radiography wide and irregular round opacity in lower right zone | 0
suspected cancer | -168
thoracoabdominal computed tomography scan performed a week ago | -168
11 cm × 9 cm × 8 cm solid mass neighboring heart | -168
surrounding atelectasis | -168
mediastinal lymphadenopathies | -168
multiple liver metastases | -168
biopsy conducted with bronchoscopy 3 days ago | -72
admitted to intensive care unit | 0
intravenous fluid hydration 200 ml/h | 0
antipotassium treatment (insulin infusion and potassium binders) | 0
allopurinol | 0
blood cultures drawn | 0
urine cultures drawn | 0
meropenem 2 g/day initiated | 0
unable to start rasburicase | 0
increases in creatinine | 0
increases in potassium | 0
increases in phosphorus | 0
consulted with nephrology department | 0
hemodialysis initiated | 0
pathology confirmed small-cell lung carcinoma | 0
patient died | 72
