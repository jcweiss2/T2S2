61 years old | 0
male | 0
hypertension | -8760
obesity | -8760
hyperlipidemia | -8760
shortness of breath | -336
cough | -336
fatigue | -336
muscle aches | -336
denies chest pain | -336
denies arm pain | -336
denies jaw pain | -336
no diabetes mellitus | -336
no cardiovascular disease | -336
no chronic lung disease | -336
no liver disease | -336
no kidney disease | -336
no tobacco use | -336
tachypneic | 0
hypoxic | 0
hypotensive | 0
tachycardic | 0
respiratory distress | 0
weak peripheral pulses | 0
cool extremities | 0
SARS-CoV-2 infection suspected | 0
sedation | 0
intubation | 0
norepinephrine | 0
vasopressin | 0
dobutamine | 0
sepsis workup | 0
septic shock workup | 0
positive SARS-CoV-2 | 0
negative other viral and bacterial pathogens | 0
elevated D-dimer | 0
elevated cardiac troponin I | 0
WBC 15.7 | 0
platelet 151 | 0
hemoglobin 13.6 | 0
creatinine 1.16 | 0
INR 1.5 | 0
CRP 306.8 | 0
LDH 707 | 0
IL-6 23 | 0
ferritin 2831.22 | 0
CK 86 | 0
new diffuse bilateral airspace opacities | 0
pulmonary infection | 0
pulmonary embolism suspected | 0
heparin infusion | 0
anticoagulation | 0
transthoracic echocardiography | 0
normal right ventricle size | 0
mildly elevated pulmonary arterial pressure | 0
moderate global hypokinesis of the left ventricle | 0
reduced overall systolic function | 0
ejection fraction 30-35% | 0
STEMI suspected | 0
acute coronary syndrome treatment | 0
aspirin | 0
ticagrelor | 0
dual antiplatelet therapy | 0
ECG ST elevation | 0
cardiac arrest | 24
death | 24
autopsy | 24
patent coronaries | 24
no significant atherosclerotic changes | 24
no acute myocardial infarct | 24
scattered focal ischemic changes | 24
interstitial edema | 24
increased macrophages | 24
adherent organizing left atrial thrombus | 24
thromboembolism of the left pulmonary artery | 24
pulmonary vascular microthrombi | 24
pulmonary consolidation | 24
hemorrhage | 24
hyaline membrane formation | 24
D-dimer 32 563 | 0
D-dimer 2816 | 96
D-dimer 1603 | 72
troponin 7457 | 0
troponin 5852 | 24
troponin 2214 | 48
troponin 0.768 | 72
platelets 242 | 72
platelets 294 | 48
platelets 385 | 24
INR 1.2 | 24
INR 1.2 | 48
INR 1.3 | 72
ventricular tachycardia | 24
coronary angiography | 48
widely patent left and right coronary arteries | 48
no epicardial stenosis | 48
no thrombosis | 48
left ventriculography | 48
diffuse hypokinesis | 48
ejection fraction 40-45% | 48
left ventricular end-diastolic pressure 22 mm Hg | 48
steroid therapy | 24
cardiopulmonary resuscitation | 24