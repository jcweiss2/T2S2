53 years old | 0
male | 0
admitted to the hospital | 0
long-standing left renal calculi | -6720
left-side pyelolithotomy | -6720
placement of a DJS | -6720
DJS placement was not performed under fluoroscopy guidance | -6720
postoperative imaging examinations were not performed | -6720
advised for stent removal after 5 months | -6720
KUB x-ray film showed DJS was not in the right location | 0
DJS appeared to enter into the IVC | 0
transferred to the hospital | 0
moderate flank pain | 0
normal leukocytes counts | 0
normal creatinine levels | 0
increased leukocytes counts in urine | 0
increased erythrocyte counts in urine | 0
urine culture was positive with a growth of Enterococcus faecalis | 0
color Doppler flow imaging showed small mural thrombus in the IVC | 0
treatments with anticoagulants | 0
treatments with antibiotics | 0
computed tomography urography | 24
migration of the DJS into the IVC | 24
left-side hydronephrosis | 24
percutaneous nephroscope under C-arm guidance | 48
distal coil of the DJS was visualized and removed | 48
new DJS was placed | 48
location of new DJS was confirmed by radiologic imaging | 48
transferred to intensive care unit | 48
treated with continued anticoagulants | 48
treated with continued antibiotics | 48
CDFI showed no thrombus in the IVC | 360
discharged | 384
follow-up was uneventful | 384