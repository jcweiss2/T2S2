64 years old | 0
male | 0
chronic pancreatitis | -8760
pseudocysts | -8760
ascites | -8760
abdominal pain | -24
hypoxic respiratory failure | -24
hypotension | -24
septic shock | -24
infected pancreatic pseudocyst | -24
necrotizing pancreatitis | -24
thrombosis in the portal vein | -24
splenic vein thrombosis | -24
superior mesenteric vein thrombosis | -24
anticoagulation | -24
pseudocyst drainage | 0
hematemesis | 24
gastroduodenal artery pseudoaneurysm | 24
transcatheter embolization | 24
coil embolization | 24
discharged | 432
hemothorax | 2160
pneumothorax | 2160
worsening ascites | 2160
anasarca | 2160
supratherapeutic International Normalized Ratio (INR) | 2160
Fresh Frozen Plasma transfusion | 2160
cardiac arrest | 2160
cardiopulmonary resuscitation | 2160
epinephrine administration | 2160
paracentesis | 2160
portal venous hypertension | 2160
hepatic and portal vein venography | 2160
core needle liver biopsy | 2160
porto-systemic venous pressure measurement | 2160
stent dilatation of the portal vein and SMV | 2160
stent placement | 2160
partial occlusion of the SMV stent | 168
anticoagulation resumed | 168
discharged | 192
asymptomatic | 7560
free of ascites | 7560
widely patent SMV and portal vein | 7560
no ascites | 7560
hepatopetal venous flow | 7560