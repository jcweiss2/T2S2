77 years old | 0
female | 0
admitted to the hospital | 0
height 148.5 cm | 0
weight 70 kg | 0
hypertension | -672
amlodipine | -672
carvedilol | -672
lumbar spinal stenosis | 0
L1-3 | 0
leukocyte count 7,770/ml | 0
hemoglobin level 14.1 mg/dl | 0
hematocrit 40.1% | 0
platelet count 268,000/ml | 0
central venous catheter | -24
ECG normal | 0
physical examination normal | 0
anesthesia induced | 0
propofol | 0
remifentanil | 0
rocuronium | 0
endotracheal intubation | 0
radial artery cannula | 0
cardiac output monitored | 0
stroke volume variation monitored | 0
systemic vascular resistance monitored | 0
cardiac index 2.8 L/min/m2 | 0
SVR index 2,394 dynes·sec/cm5/m2 | 0
mean arterial BP 95 mmHg | 0
heart rate 77 beats/min | 0
SVV 12% | 0
central venous pressure 13 mmHg | 0
arterial blood gas analysis | 0
pH 7.455 | 0
pCO2 32.9 mmHg | 0
pO2 203.7 mmHg | 0
hematocrit ratio 34% | 0
mean arterial BP decreased to 56 mmHg | 0.75
phenylephrine 50 µg | 0.75
mean arterial BP increased to 123 mmHg | 0.75
nicardipine 500 µg | 0.75
mean arterial BP decreased to 47-59 mmHg | 0.75
SVV 15% | 0.75
cardiac index 2.7-3.3 L/min/m2 | 0.75
SVRI 1,079-1,242 dynes·sec/cm5/m2 | 0.75
phenylephrine repeated | 0.75
packed red blood cells transfused | 1.5
hemoglobin level 11.0 mg/dl | 1.5
hematocrit 31.5% | 1.5
platelet count 144,000/ml | 1.5
norepinephrine administered | 2
vasopressin administered | 2
sugammadex 140 mg | 3
spontaneous respiration restored | 3
endotracheal tube removed | 3
transferred to PACU | 3
BP 82/64 mmHg | 3
heart rate 78 beats/min | 3
peripheral oxygen saturation 100% | 3
vasopressin initiated | 3.5
BP increased to 104/64 mmHg | 3.5
BP decreased to 82/57 mmHg | 3.75
ECG normal | 4
transthoracic echocardiography normal | 4
methylene blue administered | 4.5
BP increased to 112/66 mmHg | 4.5
vomiting | 4.5
methylene blue discontinued | 4.5
total dose of methylene blue 26 mg | 4.5
systolic BP remained above 110 mmHg | 5
norepinephrine and vasopressin tapered and stopped | 24
transferred to general ward | 48
discharged | 384