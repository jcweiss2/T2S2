60 years old | 0
male | 0
hypertension | 0
admitted to the hospital | 0
left eye swelling | -168
left eye pain | -168
left eye erythema | -168
circulatory shock | 0
sepsis | 0
intravenous antibiotics | 0
vancomycin | 0
gentamycin | 0
meropenem | 0
clindamycin | 0
fluid resuscitation | 0
oxygen supplementation | 0
diffuse left orbital cellulitis | 0
no intraorbital collection | 0
inflammatory picture | 0
respiratory compromise | 0
haemodynamic instability | 0
intubation | 0
ventilatory support | 0
vasopressor treatment | 0
multiorgan failure | 0
intravenous immunoglobulin | 0
left periorbital swelling | 0
necrosis of the upper eyelid | 0
suspected abscess of the lower eyelid | 0
debridement | 0
intra-operative findings of necrotizing fasciitis | 0
intensive care unit admission | 0
septic shock | 0
multiorgan failure management | 0
respiratory support | 0
vasopressors | 0
inotropes | 0
renal replacement therapy | 0
acute kidney injury | 0
antibiotic change | 0
ceftriaxone | 0
linezolid | 0
beta-haemolytic group A streptococcus | 0
Staphylococcus aureus | 0
persistent soft tissue swelling | 168
discharge | 456
wound healing | 2160
no visual deficit | 2160
awaiting reconstructive surgery | 2160
ectropion | 2160
