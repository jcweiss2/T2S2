46 years old | 0
    man | 0
    chronic bilateral hip and leg pain | 0
    left sacral fracture | 0
    sacro-iliac joint separation | 0
    tingling sensation | 0
    lancinating pain bilaterally in the hip and both legs | 0
    VAS 8 mm | 0
    motor weakness of the lower extremities | 0
    moderate sensory weakness of the lower extremities | 0
    left lumbosacral plexopathy | 0
    right chronic L5-S1 radiculopathy | 0
    acetaminophen/tramadol tablet 3 times a day | 0
    imipramine 25 mg 3 times a day | 0
    divalproate 500 mg twice a day | 0
    pregabalin 75 mg twice a day | 0
    lumbar sympathetic ganglion block | 0
    pain did not improve | 0
    Pethidine HCl 75 mg administered intravenously 4 or 5 times a day | 0
    VAS 4-8 mm | 0
    patient-controlled continuous epidural morphine infusion | 0
    preservative free morphine at a concentration of 0.28 mg/ml | 0
    basal rate of 0.5 ml/h | 0
    on-demand bolus dose of 4.0 ml | 0
    lock out interval of 30 minutes | 0
    no significant adverse events | 0
    20% pain reduction | 0
    no further improvement in pain intensity | 0
    increased basal rate up to 1.0 ml/h | 0
    considered neuromodulation | 0
    implantation of an intrathecal morphine pump | 0
    epidural PCA stopped | 0
    intrathecal morphine administration 0.3 mg | 0
    60% pain reduction | 1
    respiratory rate 17/min | 1
    pain recurred | 8
    VAS 7 | 8
    Tramadol 50 mg injected | 15
    epidural PCA restarted | 15
    dysarthria | 15
    drowsiness | 15
    no response to painful stimulation | 21
    epidural PCA stopped | 21
    unresponsive | 25
    respiratory rate 15/min | 25
    blood pressure 88/54 mmHg | 25
    oxygen saturation 69-71% | 25
    oxygen mask with reservoir bag placed | 25
    transferred to intensive care unit | 25
    Naloxone 0.4 mg administered intravenously | 25
    chest radiograph multifocal patchy consolidation | 25
    aspiration pneumonia | 25
    antibiotic therapy | 25
    ventilation care | 25
    blood gas within normal range | 72
    mentally alert | 72
    extubation | 72
    chest radiograph improved | 72
    discharged | 72
    VAS score 7 | 72