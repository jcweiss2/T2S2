23 years old | 0
male | 0
medical student | 0
disease relapse | -3456
early T-cell precursor lymphoblastic leukemia | -3456
allogenic stem cell transplantation (SCT) | -3456
re-induction therapy | -336
local radiotherapy | -336
systemic chemotherapy | -336
nelarabine | -336
triple intrathecal chemotherapy | -336
complete disease remission | -336
consolidation chemotherapy | -168
second allogenic SCT | 0
Graft-versus-host disease (GvHD) prophylaxis | 0
cyclosporine | 0
methotrexate | 0
mild oral mucositis | 120
headache | 240
moderate abdominal discomfort | 240
elevated C-reactive protein (CRP) | 240
elevated potassium levels | 240
cyclosporine dosage reduced | 240
initial improvement of symptoms | 240
recurrent hyperpotassemia | 288
SPS orally | 288
progressive abdominal pain | 288
fever | 288
body temperature 38.5°C | 288
heart rate 91 beats per minute | 288
blood pressure 126/80 mmHg | 288
peripheral oxygen saturation levels 95% | 288
bloated abdomen | 288
no signs of peritonitis | 288
low white blood cell count | 288
low neutrophils | 288
elevated CRP levels | 288
thoracoabdominal computed tomography (CT) scan | 288
thickened gastric wall | 288
gastric pneumatosis (GP) | 288
air in the hepatic portal vein system | 288
upper GI endoscopy | 300
generalized mucosal erythema | 300
intramucosal bleeding | 300
necrosis | 300
exploratory laparotomy | 312
necrosis of the gastric wall | 312
total gastrectomy | 312
end-to-side esophago-jejunal stapler anastomosis | 312
postoperative stay on the intensive care unit | 312
pain-control | 312
transferred back to the isolation ward | 312
recovered slowly | 312
total parenteral nutrition | 312
antibiotic therapy | 312
histopathology | 312
resected stomach | 312
GP | 312
circumscribed ischemic transmural necrosis | 312
purulent peritonitis | 312
kayexalate crystals | 312
no evidence of GvHD | 312
no signs of Helicobacter pylori infection | 312
vital resection margins | 312
upper GI X-ray series | 432
normal passage through the esophago-jejunostomy | 432
no signs of leakage | 432
fully recovered | 720
discharged | 720