27 years old | 0
    male | 0
    fell from 4m height | 0
    U shaped metallic bar penetrated left pelvis | 0
    trajectory toward right femur through pelvic cavity | 0
    bystanders lifted patient with bar in place | 0
    EMS arrived | -75
    hemodynamically stable | -75
    severe pain | -75
    deformed right lower extremity | -75
    evaluation by EMS staff | -75
    stabilization by EMS staff | -75
    transported to tertiary hospital | -75
    airway patent | 0
    bilateral good air entry | 0
    BP 110/70 | 0
    PR 98 | 0
    RR 12 | 0
    temperature 36.9°C | 0
    oxygen saturation 99% | 0
    GCS 15 | 0
    impaling bar found penetrating left pelvis | 0
    no active external bleeding | 0
    initial evaluation in TRU | 0
    ATLS protocol followed | 0
    FAST inconclusive | 0
    right thigh deformity | 0
    distal pulses intact | 0
    rectal exam negative for blood | 0
    rectal exam negative for masses | 0
    rectal exam negative for foreign body | 0
    prophylactic antibiotic given | 0
    tetanus toxoid given | 0
    pelvic X-ray showed right femur fracture | 0
    abdominal X-ray showed right femur fracture | 0
    protruded metal bar cut | 0
    CT scan abdomen/pelvis | 0
    metallic bar entered left pelvis | 0
    no exit site | 0
    bar passed left iliac bone | 0
    comminuted fracture supra-acetabular region | 0
    hematoma | 0
    surgical emphysema | 0
    soft tissue injury extending to left psoas muscle | 0
    bar passed junction descending/sigmoid colon | 0
    contrast extravasation | 0
    large free air upper abdomen | 0
    bar traversed soft tissue behind rectus muscle | 0
    soft tissue contusions | 0
    small metal fragment anterior to right rectus muscle | 0
    exploratory laparotomy | 0
    metallic bar removed | 0
    sigmoid colon injury | 0
    minimal contamination | 0
    sigmoid colon repair with 3-0 Vicryl sutures | 0
    thorough irrigation | 0
    systematic abdominal exploration | 0
    abdomen closed | 0
    intramedullary nailing for right femur fracture | 0
    fever | 96
    tachycardia | 96
    tachypnea | 96
    desaturation | 96
    low WBC count | 96
    intubation | 96
    admitted to ICU | 96
    broad spectrum antibiotics started | 96
    chest CT scan | 96
    abdominal CT scan | 96
    CT scan unremarkable | 96
    blood culture positive for MSSA | 96
    condition improved | 120
    extubated | 120
    transferred to ward | 144
    abdominal wound infection | 192
    pus collection | 192
    pus drained | 192
    culture positive for E. coli | 192
    antibiotic changed | 192
    wound managed | 192
    wound closed | 216
    discharged home | 240
    