4 years old | 0
male | 0
unremarkable medical history | 0
unremarkable family history | 0
admitted to the emergency room | 0
malaise | -48
lethargy | -48
tachypnea | -48
sore throat | -48
abdominal pain | -48
vomiting | -48
dehydration | -48
polyuria | -72
polydipsia | -72
weight loss | -72
afebrile | 0
tachypneic | 0
Kussmaul respirations | 0
heart rate 156 beats per minute | 0
blood pressure 90/55 mm Hg | 0
light drowsiness | 0
no jugular distension | 0
diffuse rhonchi in all lung areas | 0
diabetic ketoacidosis | 0
plasma glucose level 29.8 mmol/L | 0
pH 6.788 | 0
pO2 5.20 kPa | 0
pCO2 4.43 kPa | 0
bicarbonate 4.7 mmol/L | 0
sodium 135 mmol/L | 0
potassium 5.1 mmol/L | 0
glucosuria | 0
ketonuria | 0
insulin infusion | 0
intravenous saline | 0
potassium replacement | 0
symptomatic respiratory treatment | 0
hypotension | 0
volume expansion | 0
vasopressors | 0
inotropes | 0
severe dyspnea | 2
increased tachypnea | 2
restlessness | 2
cyanosis | 2
diffuse crackles and rhonchi in all lung areas | 2
hypoxemia | 2
bilateral severe diffuse infiltrates | 2
no cardiomegaly | 2
acute respiratory failure | 2
ARDS | 2
oxygen by facemask | 2
endotracheal intubation | 4
mechanical ventilation | 4
throat culture positive for group A beta-hemolytic streptococci | 4
intravenous co-amoxiclav | 4
intubated | 0
mechanically ventilated | 0
sedated | 0
diffusely edematous | 0
leukocyte count 18.3 | 0
differential of 67 neutrophils | 0
differential of 25 lymphocytes | 0
differential of 7 monocytes | 0
differential of 1 eosinophil | 0
prothrombin time normal | 0
platelet count normal | 0
troponin T level normal | 0
liver function tests normal | 0
levels of serum and urine amylase normal | 0
glucosuria | 0
cultures of tracheal tube negative | 0
cultures of urine negative | 0
cultures of blood negative | 0
electrocardiography pattern normal | 0
bilateral areas of patchy abnormalities | 0
mixed ground-glass appearance and consolidation | 0
no cardiomegaly | 0
no mediastinal lymphadenopathy | 0
antibiotics continued for 10 days | 0
subcutaneous injections of regular insulin | 24
euglycemia | 24
no ketonuria | 24
weaned from ventilator | 72
euglycemic | 72
no ketonuria | 72
respiratory symptoms cleared | 168
chest x-ray improved | 168
discharged | 168