50 years old | 0
male | 0
admitted to the emergency department | 0
cough | -168
phlegm | -168
sore throat | -168
fever | -96
shortness of breath | -96
chest tightness | -96
dizziness | -96
no chills | -96
no chest pain | -96
no hemoptysis | -96
no abdominal pain | -96
no diarrhea | -96
white blood cell count 8.98×10^9/L | -96
neutrophil ratio 90.7% | -96
hs-CRP 185.61 mg/L | -96
PCT 7.93 ng/mL | -96
IL-6 239.3 pg/mL | -96
CPK 2554 U/L | -96
CPK-MB 10.62 µg/L | -96
LDH 1673 U/L | -96
GOP 513.4 U/L | -96
GPT 183.1 U/L | -96
chest CT right lower lung infection | -96
enlarged right thyroid lobe | -96
black loose stools | -96
increased urination frequency | -96
urgency urination | -96
no weight changes | -96
history of thyroid enlargement | -240
Chinese medicine intake | -240
black stools history | -240
denied poultry exposure | 0
body temperature 36.6°C | 0
pulse 107 beats/min | 0
breathing 32/min | 0
blood pressure 132/97 mmHg | 0
oxygen saturation 85% | 0
FiO2 50% | 0
alert | 0
reactive pupils | 0
enlarged thyroid class II | 0
pharyngeal swelling | 0
no tonsillar swelling | 0
coarse breath sounds | 0
wet rales right lower lung | 0
heart rate 107 beats/min | 0
normal heart rhythm | 0
no murmurs | 0
no abdominal tenderness | 0
no rebound tenderness | 0
no leg edema | 0
sepsis diagnosis | 0
severe pneumonia diagnosis | 0
multiple organ dysfunction | 0
respiratory failure | 0
myocardial damage | 0
impaired liver function | 0
gastrointestinal bleeding | 0
hypokalemia | 0
hyponatremia | 0
hypochloremia | 0
blood pH 7.479 | 0
pCO2 29.3 mmHg | 0
pO2 51 mmHg | 0
base excess -2 mmol/L | 0
platelet count 94×10^9/L | 0
neutrophil ratio 92% | 0
BUN 84 µmol/L | 0
Cr 84 µmol/L | 0
hs-CRP 219.85 mg/L | 0
PCT 12.96 ng/mL | 0
CPK 18821 U/L | 0
LDH 1622 U/L | 0
GOP 395.5 U/L | 0
GPT 181.4 U/L | 0
urinary protein 3.0 g/L | 0
red blood cells 200/µL | 0
normal coagulation | 0
negative hepatitis B | 0
negative syphilis | 0
negative HIV | 0
negative hepatitis C | 0
negative influenza antigen | 0
negative bird flu | 0
negative bacterial smears | 0
negative fungal smears | 0
negative acid-fast smears | 0
negative sputum smear | 0
negative blood cultures | 0
urine culture <100 CFU/mL | 0
negative Mycoplasma antibody | 0
negative Streptococcus pneumoniae antigen | 0
negative GM test | 0
negative G test | 0
negative cryptococcal antigen | 0
negative tuberculosis immunoassay | 0
rubella IgG 34.9 IU/mL | 0
CMV IgG 189.3 AU/mL | 0
negative TORCH IgM | 0
negative CMV nucleic acid | 0
negative fecal occult blood | 0
chest radiograph right lung infection | 0
right pleural effusion | 0
endotracheal intubation | 17
mechanical ventilation | 17
imipenem/cilastatin | 17
linezolid | 17
oseltamivir | 17
methylprednisolone 80 mg | 17
worsening condition | 17
chest radiograph aggravation | 24
decreased radiolucency right lung | 24
patchy shadows left lung | 24
acute renal failure | 48
BUN 13.43 mmol/L | 48
Cr 210 µmol/L | 48
PCT 35.57 ng/mL | 48
lactic acid 2.13 mmol/L | 48
IL-6 2048 pg/mL | 48
CPK 13371 U/L | 48
CK-MB 160 U/L | 48
bronchoscopy | 72
BALF NGS | 72
blood NGS | 72
C. psittaci detection BALF | 120
C. psittaci detection blood | 120
chest CT aggregated infection | 120
increased consolidation | 120
meropenem | 120
doxycycline | 120
ceftazidime | 240
doxycycline continued | 240
weaned off ventilation | 264
tracheal extubation | 264
oral doxycycline | 264
chest CT improvement | 336
pleural effusion | 336
BUN 4.3 mmol/L | 336
Cr 47 µmol/L | 336
PCT 0.15 ng/mL | 336
lactic acid 1.7 mmol/L | 336
IL-6 9.1 pg/mL | 336
CPK 99 U/L | 336
CK-MB 22.4 U/L | 336
GOP 28 U/L | 336
GPT 48 U/L | 336
discharge | 504
diagnosis severe pneumonia | 504
ARDS | 504
sepsis | 504
multiple organ dysfunction | 504
euthyroid sick syndrome | 504
follow-up refused | 504
good physical condition | 504
