71 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
admitted to the hospital | 0 | 0 | Factual
unconscious state | 0 | 0 | Factual
history of hypertension | -720 | 0 | Factual
history of ischaemic heart disease | -720 | 0 | Factual
history of peripheral vascular disease | -720 | 0 | Factual
stroke | 0 | 0 | Factual
head computed tomographic scan | 0 | 0 | Factual
condition deteriorated rapidly | 48 | 48 | Factual
inotropic support | 48 | 48 | Factual
septic shock | 48 | 48 | Factual
elevated levels of inflammatory markers | 48 | 48 | Factual
erythrocyte sedimentation rate | 48 | 48 | Factual
C-reactive protein | 48 | 48 | Factual
blood culture | 48 | 48 | Factual
yeast in blood culture | 48 | 48 | Factual
caspofungin administered | 48 | 48 | Factual
died | 72 | 72 | Factual
Lodderomyces elongisporus identified | 72 | 72 | Factual
VITEK 2 yeast identification system | 72 | 72 | Factual
CHROMagar Candida | 72 | 72 | Factual
acetate ascospore agar | 72 | 72 | Factual
internally transcribed spacer region of ribosomal DNA sequenced | 72 | 72 | Factual
antifungal susceptibility determined | 72 | 72 | Factual
Etest | 72 | 72 | Factual
RPMI 1640 medium | 72 | 72 | Factual
glucose | 72 | 72 | Factual
amphotericin B | 72 | 72 | Factual
fluconazole | 72 | 72 | Factual
voriconazole | 72 | 72 | Factual
posaconazole | 72 | 72 | Factual
itraconazole | 72 | 72 | Factual
flucytosine | 72 | 72 | Factual
caspofungin | 72 | 72 | Factual
micafungin | 72 | 72 | Factual
no apparent risk factors | 0 | 0 | Factual
no antibiotics | 0 | 0 | Factual
no central lines | 0 | 0 | Factual
hospitalized earlier for lower limb ischaemia | -336 | -336 | Factual
discharged 2 weeks before | -336 | -336 | Factual
possibility of inoculation of the yeast from the skin | 0 | 72 | Possible
possibility of translocation from the gastrointestinal tract | 0 | 72 | Possible
Lodderomyces elongisporus is a recognized bloodstream pathogen | 0 | 0 | Factual
little is known about its virulence attributes | 0 | 0 | Factual
little is known about its environmental niche | 0 | 0 | Factual
global prevalence | 0 | 0 | Factual
isolated from patients in distant geographic regions | 0 | 0 | Factual
four patients died | 0 | 72 | Factual
six patients were treated with antifungal drugs | 0 | 72 | Factual
use of echinocandins | 48 | 72 | Factual
caspofungin | 48 | 72 | Factual
micafungin | 48 | 72 | Factual
antifungal susceptibility of L. elongisporus is scanty | 0 | 0 | Factual
no susceptibility breakpoints are available | 0 | 0 | Factual
in vitro MIC values for antifungal drugs | 72 | 72 | Factual
within the susceptible range | 72 | 72 | Factual
echinocandins have lower in vitro activity | 0 | 0 | Factual
against C. parapsilosis complex members | 0 | 0 | Factual
Infectious Disease Society of America guidelines | 0 | 0 | Factual
favour therapeutic use of echinocandins | 0 | 0 | Factual
for the treatment of candidaemia caused by C. parapsilosis | 0 | 0 | Factual
uncommon yeast pathogens are often misidentified | 0 | 0 | Factual
due to limitations of commercial yeast identification systems | 0 | 0 | Factual
VITEK 2 | 0 | 0 | Factual
does not distinguish C. parapsilosis, C. orthopsilosis, C. metapsilosis and L. elongisporus | 0 | 0 | Factual
multiplex PCR assay | 0 | 0 | Factual
simultaneously detected C. parapsilosis, C. orthopsilosis, C. metapsilosis and L. elongisporus | 0 | 0 | Factual
matrix-assisted laser desorption/ionization time-of-flight mass spectrometry | 0 | 0 | Factual
used for the identification of L. elongisporus | 0 | 0 | Factual
rare yeast species often exhibit reduced susceptibility | 0 | 0 | Factual
to one or more commonly used antifungal agents | 0 | 0 | Factual
prolonged survival of seriously ill patients | 0 | 0 | Factual
administration of multiple broad-spectrum antibiotics | 0 | 0 | Factual
dependence on life support systems | 0 | 0 | Factual
extended use of intravascular catheters | 0 | 0 | Factual
selection pressure created by prophylactic and therapeutic use of antifungal agents | 0 | 0 | Factual
resulting in increased colonization and invasive infection | 0 | 0 | Factual
delay in accurate identification | 0 | 0 | Factual
lack of experience in the management of rare yeast infections | 0 | 0 | Factual
diagnostic and therapeutic challenges | 0 | 0 | Factual
consequently higher mortality rates | 0 | 0 | Factual