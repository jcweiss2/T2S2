51 years old | 0
    woman | 0
    general convulsions | -24
    found at home lying under a pendulum clock | -24
    bolus of diazepam 20 mg | -24
    partial vigilance restored | -24
    carried to the emergency room | -24
    hypertension | -8760
    diabetes mellitus | -8760
    personality disorder | -8760
    alcohol abuse | -8760
    normal vital signs | 0
    normal physical examination | 0
    laboratory exams | 0
    tests for alcohol and drugs negative | 0
    whole-body CT scan negative for fractures or intracranial haemorrhage | 0
    pyometra due to extraneous body inside uterine cavity | 0
    focal epileptic activity in left fronto-parietal portion of brain | 0
    infusion of levetiracetam | 0
    infusion of valproate | 0
    ineffective in controlling incoming attacks | 0
    continuous administration of propofol | 0
    continuous administration of phenytoin 500 mg in 24 h | 0
    intubation | 0
    admission to ICU | 0
    endoscopic removal of extraneous body | 24
    antibiotic treatment with clindamycin | 24
    antibiotic treatment with gentamicin | 24
    hospitalization in ICU prolonged for over 5 days | 168
    progressive worsening of laboratory parameters | 168
    progressive worsening of hemodynamic parameters | 168
    hypotension | 168
    suggesting septic shock | 168
    escalation of antibiotic therapy with anidulafungin | 168
    escalation of antibiotic therapy with ceftriaxone | 168
    norepinephrine infusion 1 µg/kg/min | 168
    epinephrine infusion 1 µg/kg/min | 168
    sustained ventricular tachycardia | 180
    resolved with amiodarone 300 mg bolus | 180
    ventricular tachycardia relapsed pulseless | 180
    DC-shock | 180
    complete recovery of sinus rhythm | 180
    electrocardiogram showing diffuse ST-segment elevation | 185
    echocardiogram showing severe reduction of left ventricular function | 185
    akinesia of apex and periapical segments | 185
    apical ballooning | 185
    coronary angiography performed | 185
    coronary tree normal except mild stenosis of mid-left anterior descending artery | 185
    suggesting Tako-Tsubo syndrome | 185
    mild troponin elevation | 185
    multiple aetiologies hypothesized for TTC | 185
    substitution of phenytoin with levetiracetam | 185
    vasopressors stopped | 185
    single antiplatelet therapy with aspirin | 185
    beta-blockers started | 185
    ramipril re-introduced | 185
    extubated | 216
    discharged from ICU | 216
    progressive resolution of ST-segment elevation | 216
    recovery of left ventricular function | 216
    echocardiogram at discharge showing EF 60% | 600
    therapy with aspirin | 600
    therapy with ramipril | 600
    therapy with beta-blockers | 600
    asymptomatic at 6 months follow-up | 4320
    no further cardiovascular event | 4320
