48 years old | 0
male | 0
testicular cancer | -672
right testicular seminoma | -672
pT4 | -672
liver metastases | -672
RPLN metastasis | -672
RPLN metastasis invaded the third portion of the duodenum | -672
hCG level of 24 IU/L | -672
LDH at 1060 IU/L | -672
normal alfa-fetoprotein | -672
BEP regimen | -672
bleomycin | -672
etoposide | -672
cisplatin | -672
cisplatin dose reduced to 90% | -672
four cycles of BEP | -672
BEP regimen completed | -168
hCG normalized | -168
LDH normalized | -168
contrast-enhanced CT | -168
PET-CT | -168
disappearance of liver metastases | -168
RPLN mass remained | -168
positive 18F-FDG uptake | -168
referred to hospital | -84
RPLND considered | -84
repeat PET-CT | -84
increasing 18F-FDG uptake | -84
new uptake in right iliac lymph node metastases | -84
salvage chemotherapy | -84
paclitaxel | -84
ifosfamide | -84
TIP treatment | -84
no severe adverse effects | -84
CT after two courses of TIP | -42
RPLN metastasis did not respond to chemotherapy | -42
adverse effect of two additional courses of TIP | -42
sudden-onset hematochezia | 0
hypovolemic shock | 0
hemoglobin 4.7 g/dL | 0
neutrophil count 4.8 × 10^9/L | 0
platelet count 4.9 × 10^9/L | 0
CT depicted dilated bowel loop | 0
massive clot | 0
direct extravasation of contrast from aorta into duodenum | 0
RPLN mass remained without decrease in size | 0
endoscopic therapy considered impossible | 0
angioembolization attempted | 0
emergent angiography | 0
PADF confirmed | 0
endovascular stent graft deployed | 0
control angiography | 0
minimal residual hemorrhage | 0
extensive fluid infusion | 0
blood transfusion | 0
sepsis | 24
DIC | 24
MOF | 24
definitive surgical repair awaited | 24
massive bleeding recurred | 432
patient died | 432
septic shock | 432
uncontrolled bleeding | 432