62 years old | 0
woman | 0
alcohol abuse | -72
dental pain | -72
facial swelling | -72
altered mental status | -72
admitted to the emergency department | 0
Glasgow Coma Scale 13 | 0
disoriented to time | 0
disoriented to place |7
febrile | 0
temperature 40° Celsius | 0
heart rate 160 beats per minute | 0
hypertension | 0
family history of seizure disorder | 0
daily alcohol intake | 0
pupils 1 mm | 0
minimally reactive to light | 0
no afferent pupillary defect | 0
visual acuity hand motion | 0
orthotropic in primary gaze | 0
full ocular motility | 0
intraocular pressure 19 mm Hg right | 0
intraocular pressure 14 mm Hg left | 0
right periorbital edema | 0
right temporal edema | 0
right periorbital erythema | 0
right temporal erythema | 0
inferior chemosis right conjunctiva | 0
no conjunctival erythema | 0
unremarkable fundus examination | 0
septic shock | 0
serum anion gap 23 mEq/L | 0
lactic acid 4.8 mmol/L | 0
white blood cell count 15,000/mm3 | 0
intravenous vancomycin | 0
intravenous piperacillin/tazobactam | 0
intravenous metronidazole | 0
unremarkable urinalysis | 0
chest radiograph right upper lung opacity | 0
chest radiograph basilar opacities | 0
CT chest bilateral lung masses | 0
CT chest nodules with feeding vessel sign | 0
CT face multi-fascial space abscesses | 0
CT face phlegmon | 0
CT face gas extending to right lateral supraorbital soft tissues | 0
thrombophlebitic right retromandibular vein | 0
thrombophlebitic right superior temporal vein | 0
periorbital cellulitis | 0
thrombophlebitis right infraorbital facial vein | 0
thrombophlebitis right internal jugular vein | 0
unremarkable CT head | 0
transthoracic echocardiogram | 0
mild to moderate aortic regurgitation | 0
small pericardial effusion | 0
no valvular vegetation | 0
no intracardiac abscess | 0
incision and drainage facial abscesses | 72
extraction of five carious teeth | 72
Streptococcus constellatus identified | 72
negative tracheal aspirate | 72
negative urine cultures | 72
vancomycin discontinued | 72
clindamycin discontinued | 72
piperacillin/tazobactam discontinued | 72
ampicillin/sulbactam started | 72
anticoagulation considered | 72
anticoagulation held | 72
eradication of bacteremia | 72
transferred out of ICU | 168
binocular diplopia | 168
right incomitant esotropia | 168
-4 abduction defect | 168
lateral rectus paralysis | 168
right sixth nerve palsy | 168
intact cranial nerve function | 168
intact extraocular movements | 168
no nystagmus | 168
intraocular pressure 16 mm Hg | 168
visual acuity 20/30 bilaterally | 168
mild chemosis | 168
improved chemosis from admission | 168
no conjunctival erythema | 168
CT angiogram hypoenhancement cavernous sinuses | 168
persistent multifascial abscesses | 168
repeat incision and drainage | 168
anticoagulation considered again | 168
anticoagulation avoided due to gastrointestinal bleed | 168
another incision and drainage | 168
discharged | 168
switched to ertapenem | 168
no improvement of sixth nerve palsy | 1008
