67 years old | 0
male | 0
admitted to the intensive care unit | 0
suspected sepsis | 0
isolation of alpha-hemolytic Streptococcus pneumoniae from blood culture | 0
Gram stain revealing lanceolate diplococci | 0
positive capsule staining by India ink | 0
optochin resistance | 0
bile solubility | 0
inulin fermentation | 0
identification by VITEK II | 0
identification by MALDI-TOF | 0
detection of lytA gene | 0
detection of ply gene | 0
gene sequencing showing synonymous single nucleotide polymorphism in lytA gene | 0
treatment with ceftriaxone | 0
discharge after complete recovery | 24
