18 years old | 0
male | 0
splenectomy | -43
idiopathic thrombocytopenic purpura | -43
menometrorhagia | -43
PPV23 | -43
idiopathic thrombocytopenic purpura treatment | -43
menometrorhagia treatment | -43
vaccination with PPV23 | -43
splenectomy due to idiopathic thrombocytopenic purpura | -43
general body malaise | -2
diarrhea | -2
vomiting | -2
influenza-like symptoms | -2
increasingly more confused | 0
fever | 0
hypotension | 0
bradycardia | 0
tachypnea | 0
decreased oxygen saturation | 0
cyanosis of the lips and distal extremities | 0
sepsis | 0
volume therapy | 0
broad-spectrum antimicrobial therapy | 0
hydrocortisone | 0
white blood cell count | 0
neutrophils | 0
hemoglobin | 0
thrombocytes | 0
C-reactive protein | 0
P-lactate | 0
aB-P-O2 | 0
aB-P-CO2 | 0
aB-pH | 0
Streptococcus pneumococcal urinary antigen test positive | 0
chest x-ray | 0
disseminated intravascular coagulation | 24
microthrombi in the hands and feet | 24
blood cultures showed growth of S. pneumoniae | 24
antimicrobial treatment changed to penicillin G | 24
modest hypokinesia of the apical part of the left ventricle | 48
ejection fraction of 45% | 48
endocarditis dismissed | 48
necrosis of the fingertips and toes | 48
renal insufficiency | 48
hemodialysis | 48
antibiotic therapy altered to ceftriaxone | 48
leucocytes and CRP decreased | 96
fever dissolved | 96
tracheal secret for culture had been obtained | 96
culture was negative | 96
transferred from the ICU to the medical department | 144
antibiotics were stopped | 144
serological analysis of the pneumococcal isolate | 144
serotype 12F | 144
afebrile with fluctuating CRP | 155
condition improved clinically | 155
discharged with oral dicloxacillin | 155
raised leucocytes and CRP | 155
site of current infection suspected to be the necrotic tissue | 155
wound cultures had shown Staphylococcus aureus and haemolytic streptococci group C/G | 155
new TTE was unchanged | 155
necrotic fingers and toes were amputated | 168
readmitted with severe sepsis | 213
sepsis regimen and ceftriaxone therapy | 213
transesophageal echocardiography revealed endocarditis | 213
blood cultures showed growth of S. pneumoniae | 213
antimicrobial treatment altered to penicillin G | 213
penicillin G for 4 weeks | 217
recovered | 217
serological tests of the pneumococcal capsule polysaccharides | 217
serotype 12F | 217
serological tests of the pneumococcal capsule polysaccharides | 217
serotype 12F | 217
serological tests of the pneumococcal capsule polysaccharides | 217
serotype 12F | 217
investigated whether the patient was able to respond to serotype 12F with antibodies | 217
confirmed a 12F-antibody response | 217
antibody response was not great enough to avoid IPD | 217