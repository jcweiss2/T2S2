54 years old | 0
lady | 0
HIV infection | -175200
pain over the right hip | 0
inability to bear weight on the right lower limb | 0
trivial fall | 0
first-line ART | -52560
TDF 300 mg | -52560
lamivudine 300 mg | -52560
efavirenz 600 mg | -52560
tenderness over the right hip | 0
shortening of the right lower limb | 0
restricted range of motion | 0
fractured neck of the right femur | 0
admitted | 0
planned for hemiarthroplasty | 0
azotemia | 0
hypokalemia | 0
anemia | 0
glycosuria | 0
proteinuria | 0
raised serum alkaline phosphatase level | 0
normal anion gap metabolic acidosis | 0
glucose 3+ | 0
protein 1+ | 0
few red blood cells | 0
oral potassium supplementation | 0
ART modified to abacavir 600 mg | 0
lamivudine 150 mg OD | 0
efavirenz 600 mg OD | 0
diagnosis of renal Fanconi syndrome | 0
hypophosphatemia | 0
hyperchloremic metabolic acidosis | 0
gross dilatation of the right kidney's pelvicalyceal system | 0
multiple calculi involving both the kidneys | 0
four calculi in the right kidney's lower polar region | 0
6-mm calculus in the proximal right ureter | 0
upstream hydroureteronephrosis | 0
3-mm calculus in the lower polar calyx of the right kidney | 0
cystopanendoscopy | 0
right double "J" stenting | 0
tachycardia | 72
tachypnea | 72
hypotension | 72
pulmonary thromboembolism | 72
unfractionated heparin | 72
neutrophilic leucocytosis | 78
worsening azotemia | 78
severe metabolic acidosis | 78
urine culture grew Escherichia coli | 78
urine culture grew Enterobacter aerogenes | 78
postoperative urinary tract infection | 78
culture-sensitive injectable antibiotics | 78
bicarbonate infusion | 78
serum creatinine improved to 1.4 mg/dL | 96
discharged | 96
no orthopedic intervention | 96
advice to follow up after 1 month | 96
