74 years old | 0
male | 0
hypertension | -672
insulin-dependent diabetes mellitus type 2 | -672
diabetic retinopathy | -672
weight loss | -168
iron deficiency anemia | -168
tumor in the colon ascendens | -168
liver metastases | -168
right hemicolectomy | -24
low-grade pT3cN0 adenocarcinoma | -24
absence of metastases in 24 excised lymph nodes | -24
lymphovascular growth | -24
no vascular or perineural growth | -24
activated BRAF mutation in exon 15 (V600E) | -24
loss of expression of MLH1 and PMS2 | -24
mismatch repair-deficient (MMR-D)/microsatellite-instable (MSI) tumor | -24
initiated therapy with pembrolizumab | 0
symptoms of a cold | 7
leukocytosis | 7
slight increase in C-reactive protein | 7
dry coughing | 22
no fever | 22
increase in AST and ALT | 22
ICI-induced hepatitis grade 2 | 22
initiated prednisolone therapy | 22
second dose of pembrolizumab not given | 22
dyspnea | 29
elevation of troponin T | 29
septal hypokinesia | 29
somnolence | 29
difficulty walking | 29
dysarthria | 30
hoarseness | 30
pain in neck and right leg | 30
difficulty raising right leg | 30
increased dose of prednisolone | 30
computed tomography did not show signs of stroke | 30
increased creatine kinase and myoglobin levels | 30
ICI-induced myositis suspected | 30
antibodies against acetylcholine receptor and titin present | 30
albumin present in cerebrospinal fluid | 30
unable to sit up | 34
severe dysarthria and dysphagia | 34
absent reflexes in biceps, brachioradialis, triceps, and patellar and Achilles tendons | 34
transferred to intensive care unit | 34
intubated | 35
given methylprednisolone | 35
given intravenous immunoglobulins | 35
given infliximab | 37
felt better and had better muscle strength in hands | 38
developed carbon dioxide retention | 39
needed noninvasive ventilation | 39
developed sinus bradycardia | 39
died | 39
significant stenosis of right coronary artery | 39
no fibrosis or signs of recent myocardial infarction | 39
softened tongue | 39
no surgical complication after hemicolectomy | 39
metastasis in right liver lobe | 39
pronounced inflammatory infiltration of lymphocytes, occasional plasma cells and granulocytes, and fibrosis in intercostal musculature, diaphragm, cervical musculature and tongue | 39
fibrosis in one area of heart | 39
inflammatory infiltrate in small area of heart | 39
hepatocellular cancer (HCC) in liver | 39
HCC positive for hepatocytes and negative for glypican, CDX2, CK20 and CK7 | 39
fibrosis stage 2–3 according to Batts and Ludwig in porta field | 39