42 years old | 0
male | 0
admitted to the hospital | 0
stage 1 S germ cell tumor of the mediastinum | -5040
hemorrhagic pituitary prolactinoma | -5040
left middle cerebral artery thrombotic stroke | -5040
Etoposide treatment | -168
Ifosfamide treatment | -168
Cisplatin treatment | -168
Cabergoline treatment | -168
febrile neutropenia | 0
septic shock | 0
Escherichia Coli bacteremia | 0
severe anemia | 0
low platelet count | 0
blood transfusions | 0
platelet transfusions | 0
respiratory failure | 0
mechanical ventilation | 0
blood pressure support | 0
norepinephrine treatment | 0
dobutamine treatment | 0
vasopressin treatment | 0
phenylephrine treatment | 0
methylprednisolone treatment | 0
meropenem treatment | 0
hematemesis | 480
drop in hemoglobin | 480
pantoprazole drip | 480
upper endoscopy | 480
blood clots in the fundus | 480
ulcers in the gastric antrum | 480
normal esophagus | 480
normal duodenum | 480
biopsy of an ulcer | 480
chronic active gastritis | 480
foveolar hyperplasia | 480
repeat endoscopy | 480
IV erythromycin | 480
multiple ulcers | 480
large blood clot in the fundus | 480
mesenteric angiography | 480
left gastric artery embolization | 480
exploratory laparotomy | 504
distended stomach | 504
blood filled stomach | 504
multiple deep ulcerations | 504
total gastrectomy | 504
esophagojejunostomy | 504
jejunostomy tube placement | 504
gross pathology | 504
multiple hemorrhagic deep ulcerations | 504
broad aseptate fungi | 504
angioinvasion | 504
Warthin Starry stain | 504
immunostaining | 504
negative for Helicobacter pylori | 504
negative for Cytomegalovirus | 504
hemodynamically stable | 528
off blood pressure support medications | 528
extubated | 528
sputum cultures | 528
Aspergillus fumigatus | 528
amphotericin B treatment | 528
voriconazole treatment | 528
renal failure | 528
isavuconazole treatment | 528
discharged to rehabilitation facility | 1008
posaconazole treatment | 1008
micafungin treatment | 1008
Mycotypha microspora | 504
invasive gastric mucormycosis | 504