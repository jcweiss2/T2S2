17 years old | 0  
    black | 0  
    African | 0  
    female | 0  
    admitted to the hospital | 0  
    gradual-onset bi-frontal headache | -336  
    insomnia | -336  
    subjective fevers | -336  
    restlessness | -240  
    third-person auditory hallucinations | -240  
    acute schizoaffective disorder | -240  
    psychological stressors | -240  
    death anniversary of her mother | -240  
    imminent final high-school national examinations | -240  
    documented fevers | -168  
    orofacial dyskinesias | -168  
    tongue-biting | -168  
    agitation | -168  
    neuroleptic malignant syndrome | -168  
    coma | -144  
    transferred to tertiary referral hospital | -144  
    temperature of 39°C | 0  
    tachycardia | 0  
    Glasgow Coma Scale 7/15 | 0  
    grimacing | 0  
    tongue biting | 0  
    bruxism | 0  
    hyper-salivation | 0  
    abnormal arm movements | 0  
    intubated | 0  
    mechanically ventilated | 0  
    admitted to intensive care unit | 0  
    elevated CSF pressures | 0  
    CSF white cell count 115/mm3 | 0  
    CSF lymphocytes 98% | 0  
    negative PCR for bacterial meningo-encephalitis pathogens | 0  
    negative PCR for tuberculosis meningo-encephalitis pathogens | 0  
    negative PCR for herpes meningo-encephalitis pathogens | 0  
    contrast-enhanced MRI brain scan leptomeningeal enhancement | 0  
    MRI sulcal hyperintensities | 0  
    EEG diffuse slowing | 0  
    EEG no epileptiform discharges | 0  
    treated for viral encephalitis | 0  
    stopped viral encephalitis treatment after negative PCRs | 0  
    probable NMDARE diagnosis | 0  
    intravenous methylprednisolone | 0  
    intravenous immunoglobulins | 0  
    oral levetiracetam | 0  
    tetrabenazine | 0  
    midazolam infusion | 0  
    propofol infusion | 0  
    maxillo-mandibular fixation | 0  
    serum positive for NMDA receptor antibodies | 7  
    CSF positive for NMDA receptor antibodies | 7  
    MRI pelvis no teratoma | 7  
    repeat MRI brain resolution of meningeal enhancement | 15*24  
    repeat MRI brain resolution of sulcal hyperintensities | 15*24  
    Glasgow Coma Scale 8/15 | 15*24  
    persistent dyskinesias | 15*24  
    repeated IVMP course | 15*24  
    plasma exchange | 15*24  
    weekly rituximab | 15*24  
    right brachial deep vein thrombosis | 15*24  
    treated with low-molecular weight heparin | 15*24  
    tongue maceration | 15*24  
    surgical debridement | 15*24  
    tracheostomy | 15*24  
    percutaneous endoscopic gastrostomy | 15*24  
    high-grade fevers | 21*24  
    multi-drug resistant Pseudomonas aeruginosa | 21*24  
    Klebsiella pneumoniae | 21*24  
    appropriate intravenous antibiotics | 21*24  
    carbapenems | 21*24  
    continued debridement | 21*24  
    septic shock | 30*24  
    multi-organ dysfunction | 30*24  
    death | 30*24  
    <|eot_id|>
    
