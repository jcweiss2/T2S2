40 years old | 0
female | 0
chronic alcoholic | 0
admitted to the hospital | 0
transient hypothermia-related acute pancreatitis | 0
hypothermic at 81°F | 0
warming blanket applied | 0
serum alcohol level 0.01 | 0
creatinine phosphokinase 564 | 0
blood urea nitrogen 16 | 0
creatinine 0.4 | 0
glucose 58 | 0
aspartate transaminase 188 | 0
alanine transaminase 69 | 0
alkaline phosphatase 216 | 0
TSH 1.07 | 0
prolactin 44.9 | 0
amylase 498 | 0
lipase 1,200 | 0
ammonia 26 | 0
serum carboxyhemoglobin level 2.4 | 0
magnesium 1.3 | 0
cortisol 38 | 0
β-HCG negative | 0
generalized tonic-clonic seizure | 8
intravenous lorazepam 2 mg | 8
levetiracetam 1,000 mg | 8
transient hypotension | 8
fluid challenge with 2 L normal saline | 8
vancomycin given | 8
cefepime given | 8
metronidazole given | 8
sepsis workup negative | 8
antibiotics held off | 8
sonogram showed fatty liver | 0
trace ascites | 0
CAT scan showed no radiopaque gallstones | 0
peripancreatic fluid | 0
fluid in splenic flexure of colon | 0
fluid inferior aspect of spleen | 0
pancreas symmetrically enhanced | 0
no pancreatic necrosis | 0
no hemorrhage | 0
no peripancreatic abscess | 0
no pancreatic mass | 0
low-fiber low-fat diet tolerated | 96
discharged | 96
