32 years old | 0
male | 0
admitted to the hospital | 0
bilateral lower extremities weakness | -48
inability to walk | -48
progressive bilateral lower extremities weakness | -2160
slurred speech | -336
deviation of the left eye | -336
hypothyroidism | -4320
acquired immune deficiency syndrome | -4320
CD4+ T-lymphocyte cell count <20 | -4320
plasma HIV RNA (viral load) of 206,000 | -4320
dysarthria | 0
horizontal nystagmus bilaterally | 0
dysmetria on finger-to-nose examination | 0
unsteady gait | 0
abnormal non-enhancing hyperintense T2 hypointense T1 signal extending from central cerebellar white matter | 0
superior cerebellar peduncles involvement | 0
pons involvement | 0
cerebral peduncles involvement | 0
left cortical spinal tract involvement |; 0
hypoxic | 120
hypotensive | 120
altered mental status | 120
intubated | 120
broad-spectrum antibiotics | 120
transferred to the ICU | 120
VRE peri-rectal surveillance cultures sent | 120
VRE peri-rectal surveillance cultures negative | 120
failed multiple weaning attempts | 168
percutaneous tracheostomy | 168
percutaneous endoscopic gastrostomy tube placement | 168
severe watery diarrhea | 504
C. difficile glutamate dehydrogenase positive | 504
C. difficile toxin B positive | 504
oral vancomycin started | 504
diarrhea persisted | 1344
bleeding per rectum | 1344
solid brown stool | 1344
specks old blood | 1344
no fresh blood | 1344
colonoscopy scheduled | 1344
diffuse area of severely altered vascular | 1344
congested mucosa | 1344
erythematous mucosa | 1344
friable with contact bleeding mucosa | 1344
hemorrhagic mucosa | 1344
inflamed mucosa | 1344
nodular mucosa | 1344
ulcerated mucosa | 1344
oral and rectal vancomycin with metronidazole started | 1344
blood culture no growth | 1344
urine culture no growth | 1344
tissue culture grew VRE | 1344
echocardiogram showed no vegetation | 1344
Infectious disease consulted | 1344
clinical condition improved | 1680
diarrhea resolved | 1680
discharged | 1680
