61 years old | 0
male | 0
admitted to the hospital | 0
acute onset rapidly progressive diffusely erythematous rash | -168
rash within the deep folds of his pannus | -168
rash in the intertriginous areas | -168
never had this type of rash previously | -168
rash refractory to over-the-counter topical nystatin therapy | -168
over-the-counter topical nystatin therapy | -168
initial presentation | 0
rash suspicious for candidal intertrigo | 0
erythrasma high on the differential diagnosis | 0
coral red florescence noted with woods lamp | 0
started empirically on oral erythromycin | 0
started empirically on oral fluconazole | 0
rash spread diffusely across his trunk | -72
rash spread to extremities | -72
erythematous morbilliform papules coalesced to form plaques | -72
worsening rash | -12
acutely decompensated | -12
became short of breath | -12
developed metabolic acidosis | -12
developed respiratory acidosis | -12
transfer to the intensive care unit | -12
started on BiPAP | -12
increasing somnolence | -12
intubated | -12
hypotensive | -12
not responsive to intravenous fluid resuscitation | -12
started on vasopressor support with norepinephrine | -12
developed shock liver | -12
developed acute kidney failure requiring CVVHD | -12
neutrophilic leucocytosis | 0
white blood cell 31.10× 109/L | 0
acute kidney failure | 0
creatinine of 3.06 mg/dL | 0
hyperkalaemia of 6.3 mmol/L | 0
phosphorus of 7.0 mg/dL | 0
metabolic acidosis | 0
respiratory acidosis | 0
shock liver | 0
AST of 4902 units/mL | 0
ALT of 3073 units/mL | 0
CXR normal | 0
CT chest/abdomen and pelvis no focal signs of infection | 0
blood culture negative for bacterial/fungal growth | 0
urine culture negative for bacterial/fungal growth | 0
superficial wound culture grew Streptococcus agalactiae | 0
superficial wound culture grew rare Proteus mirabilis | 0
superficial wound culture grew rare Klebsiella | 0
superficial wound culture grew coagulase-negative Staphylococcus | 0
skin biopsy showed diffuse spongiosis | 0
skin biopsy showed numerous subcorneal pustules | 0
mixed inflammatory infiltrate predominately neutrophils | 0
some associated lymphocytes | 0
diagnosis of AGEP | 0
septic shock less likely | 0
pustular psoriasis less likely | 0
TEN less likely | 0
SJS less likely | 0
abrupt onset | 0
short duration | 0
rapid improvement after drug withdrawal | 0
no evidence of arthritis | 0
no personal history of psoriasis | 0
no family history of psoriasis | 0
no mucous membrane involvement | 0
discontinued erythromycin | 0
discontinued fluconazole | 0
started on vancomycin | 0
started on meropenem | 0
started on micafungin | 0
antibiotics discontinued | 0
treated with methylprednisolone 80 mg every 8 hours for 3 days | 0
slow taper on oral steroids | 0
marked improvement in haemodynamics | 72
marked improvement in rash | 72
no longer required vasopressor agents | 72
extubated on day 3 | 72
required 4 days of CVVHD | 96
complete recovery of kidney function | 96
complete recovery of liver function | 96
maintained on oral prednisone | 96
slow taper for 2 weeks | 336
morbid obesity | 0
Chronic Obstructive Pulmonary Disease | 0
hypertension | 0
type 2 diabetes mellitus | 0
