40 years old | 0
male | 0
rheumatoid arthritis | -1920
immunosuppressive medication | -1920
prednisolone | -1920
hydroxychloroquine | -1920
paroxysmal AF | -168
palpitation | -168
atrial fibrillation ablation | 0
radiofrequency catheter ablation | 0
general anesthesia | 0
mechanical ventilation | 0
3-dimensional navigation system | 0
irrigation tip ablation catheter | 0
electrical isolation of pulmonary vein | 0
esophageal temperature monitoring | 0
intracardiac echocardiography | 0
ablation power | 0
temperature cutoff | 0
impedance cutoff | 0
radiofrequency ablation | 0
persistent retrosternal pain | 24
fentanyl-patch application | 24
morphine injections | 24
pantoprazole | 24
symptomatic AF recurrence | 72
bisoprolol | 72
flecainide | 72
discharged | 120
recurring symptomatic AF | 216
mild chest pain | 216
paroxysmal palpitation | 216
chest pain aggravation | 408
deep inspiration | 408
coughing | 408
fever | 408
severe chills | 408
leukocytosis | 408
normal sinus rhythm | 408
cardiac troponin-I | 408
C-reactive protein | 408
no cardiomegaly | 408
no pleural effusion | 408
abnormal pericardial fluid collection | 408
chest computed tomography | 408
small air bubbles in pericardial space | 408
esophageal perforation | 408
admitted to sub-intensive care unit | 408
broad-spectrum antibiotics | 408
sepsis | 480
multi-organ failure | 480
pericardial and pleural effusions | 480
large air bubbles in pericardial space | 480
esophagography | 480
contrast agent leakage into pericardial space | 480
pericardiostomy | 480
chest tubing | 480
pericardial drainage tube | 480
strict fasting | 480
fluid replacement | 480
broad-spectrum antibiotic therapy | 480
continuous drainage | 480
recovered from sepsis | 504
recovered from multi-organ failure | 504
follow-up esophagography | 624
no contrast agent leakage | 624
dietary intake restarted | 624
follow-up chest CT | 720
improving mediastinitis | 720
discharged | 1008
antiarrhythmic therapy | 1008
administration of antiarrhythmic agents stopped | 2160