32 years old | 0
male | 0
admitted to the hospital | 0
fever | -48
cough | -48
shortness of breath | -48
diarrhea | -72
exposure to father with similar symptoms | -72
no chest pain | 0
no abdominal pain | 0
no nausea | 0
no vomiting | 0
regular heart rate | 0
regular heart rhythm | 0
no murmurs | 0
no rubs | 0
no gallops | 0
no jugular venous distension | 0
lungs clear to auscultation bilaterally | 0
ecchymosis from cupping marks | 0
normotensive | 0
no tachycardia | 0
respiratory rate 18 breaths per min | 0
oxygen saturation 95% on room air | 0
unremarkable complete blood count | 0
hyper-glycemia | 0
elevated hemoglobin A1c | 0
elevated lactate dehydrogenase | 0
elevated C-reactive protein | 0
mild acidemia | 0
normal sinus rhythm | 0
no QTc prolongation | 0
peripheral patchy opacities in the lower lung zones | 0
started on IV ceftriaxone | 0
started on IV azithromycin | 0
started on IV hydroxychloroquine | 0
started on oral zinc supplementation | 0
desaturated to 79% SpO2 | 1
required 6 L/min supplemental oxygen | 1
switched to high-flow nasal cannula | 1
added IV linezolid | 1
started insulin regimen | 1
SARS-CoV-2 RNA positive | 48
influenza A nasal swab positive | 48
added oseltamivir | 48
chest computed tomography scan | 48
extensive bilateral ground-glass opacities | 48
confluent consolidation in the posterior lung bases | 48
fever spikes | 48
worsening tachypnea | 120
increased FiO2 requirement | 120
worsening PaO2/FiO2 ratio | 120
SpO2 around 87% | 120
increased respiratory rate | 120
elevated ferritin level | 120
persistently elevated LDH level | 120
normal pH | 120
normocarbia | 120
hypoxia | 120
elevated bicarbonate level | 120
intubated | 120
placed on mechanical ventilation | 120
upgraded to Intensive Care Unit | 120
given IV tocilizumab | 120
acute kidney injury | 120
anuric | 120
started hemodialysis | 120
discontinued linezolid | 120
started IV meropenem | 120
started IV lopinavir and ritonavir | 120
self-extubated | 168
transitioned to bilevel positive airway pressure | 168
transitioned to high-flow nasal cannula | 168
downgraded | 168
found to be hypoxic on the medical floor | 168
repeat chest X-ray | 168
worsening opacities | 168
placed on bilevel positive airway pressure again | 168
went into respiratory distress | 168
re-intubated | 168
placed back in the ICU | 168
died | 240