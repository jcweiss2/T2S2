25 years old | 0
male | 0
Romanian | 0
Roma community | 0
living in France | 0
admitted to the hospital | 0
fever | -72
diarrhea | -72
conjunctivitis | -72
no history of medical or surgical disease | 0
no treatment upon admission | 0
smoked 5 cigarettes per day | 0
no risks of sexually transmitted diseases | 0
fever at 38.5°C | 0
tachycardia at 125 beats per minute | 0
sweat | 0
submandibular centimetric lymphadenopathies | 0
Koplik's spots | 0
bilateral conjunctivitis | 0
erythematous extending facial eruption | 0
diarrhea without signs of dehydration | 0
stable blood pressure at 129/68 mm Hg | 0
normal pulmonary auscultation | 0
normal neurological examination | 0
hyponatremia at 126 mmol/L | 0
hypokalemia at 3.33 mmol/L | 0
mild acute renal insufficiency | 0
elevated creatinine at 100 μmol/L | 0
clearance at 86 mL/min | 0
anicteric cholestasis | 0
cytolysis 3 times higher than normal | 0
inflammatory syndrome with C reactive protein at 55 mg/L | 0
normal chest X-rays | 0
bilateral pneumonia | 48
thoracic computed-tomography scanner | 48
diagnosis of measles | 48
positive immunoglobulin M in serum | 48
positive PCR in urine | 48
positive PCR in pharyngeal sample | 48
positive PCR in serum | 48
transferred to the intensive care unit | 72
multiorgan failure | 72
neurological failure | 72
hyponatremia | 72
acute measles encephalitis | 72
positive PCR for measles in the cerebrospinal fluid | 72
normal magnetic resonance imaging | 72
cardiac and respiratory failure | 72
septic shock | 72
bilateral associated wild type of Staphylococcus aureus and measles-linked pneumonia | 72
severe hepatic cytolysis | 72
fortuitously diagnosed hepatitis B | 72
treated with ophthalmic vitamin A for a corneous ulcer | 72
hypophosphoremia at 0.62 mmol/L | 72
severe vitamin A deficiency at 0.17 mg/L | 72
supplemented during hospitalization | 72
measles complicated with pneumonia | 72
acute encephalitis | 72
pancreatitis | 72
corneous ulcer | 72
associated with vitamin A deficiency | 72
treated with intravenous ribavirin | 72
treated with intramuscular vitamin A | 72
treated with ophthalmic vitamin A therapy | 72
pneumonia required initial intubation | 72
treated with antistaphylococcal agent | 72
successfully extubated at day 11 | 264
complete respiratory recovery | 264
complete neurological recovery | 264
complete cardiac recovery | 264
complete renal recovery | 264
complete ophthalmic recovery | 264
complete digestive recovery | 264
vitamin A control revealed normalization at 0.58 mg/L | 264
discharged | 480