61 years old | 0
male | 0
admitted to the intensive care unit | 0
nasal cavity rhinoscleroma | -672
unconscious | 0
Glasgow Coma Scale score of 10/15 | 0
tachycardic at 145 bpm | 0
hypotensive at 86/51 mm Hg | 0
polypneic at 32 cpm | 0
desaturated at 40% at room air | 0
desaturated at 78% under high mask concentration 15 L/mn | 0
body temperature was 38.5°C | 0
diffuse subcrackling rales | 0
ulcerative lesions of the nasal cavity | 0
ulcerative lesions of the oral cavity | 0
lactate level 3.24 | 0
PaO2/FiO2 ratio of 105 | 0
elevated levels of white blood cells to 14,600/µL | 0
C-reactive protein level elevated to 230 mg/L | 0
procalcitonin positive at 2.32 g/L | 0
lymphopenia at 180/µL | 0
anemia at 8.4 g/dL | 0
prothombin time at 51% | 0
high level of D-dimers 2.76 mg/L | 0
normal renal function | 0
normal hepatic function | 0
sinus tachycardia | 0
no conduction or repolarization disturbances | 0
bilateral infectious bronchopneumonia | 0
moderate bilateral pleurisy | 0
no signs of pulmonary embolism | 0
normal transthoracic echocardiogram | 0
diagnosed with pneumonia caused by Klebsiella rhinoscleromatis | 0
intubated | 0
given vasoactive drugs such as noradrenaline | 0
intravenous antibacterial treatment using Triaxon 2 g/d | 0
intravenous antibacterial treatment using ciprofloxacin 200 mg twice a day | 0
bacterium detected in a distal pulmonary swab | 24
bacterium detected in the blood culture | 24
organ dysfunction failure | 240
death | 240