57 years old | 0\
Hispanic | 0\
male | 0\
coronary artery disease | -3024\
myocardial infarction | -3024\
ischemic dilated cardiomyopathy | -3024\
pocket infection of his cardiac resynchronization therapy defibrillator | -48\
erythema around his left upper chest implant site | -720\
discomfort around his left upper chest implant site | -720\
edema around his left upper chest implant site | -720\
serosanguinous drainage around his left upper chest implant site | -720\
oral amoxicillin treatment | -720\
nonbacteremic | -48\
afebrile | -48\
severely reduced left ventricular systolic function | -48\
ejection fraction of 20%–25% | -48\
global hypokinesis of the left ventricle | -48\
no evidence of vegetations | -48\
leads were scarred to the lateral wall of the superior vena cava | -48\
transvenous lead extraction | 0\
cardiac resynchronization therapy defibrillator pocket capsule was dissected out | 0\
device removed | 0\
coronary sinus and right atrial leads were extracted | 0\
right ventricular lead was extracted | 0\
hypotensive | 0\
large pericardial effusion | 0\
emergency midsternotomy | 0\
bleeding was manually controlled with pressure | 0\
cardiopulmonary bypass was instituted | 0\
5-mm tear in the superior cavoatrial junction | 0\
perforation in the right atrium | 0\
oozing hematoma at the level of the innominate vein | 0\
repair with multiple 4-0 polypropylene sutures with pledgets | 0\
right ventricular lead was capped and abandoned | 0\
intra-aortic balloon pump was placed | 0\
hemodynamic instability | 0\
multiple blood transfusions | 0\
coagulopathy | 0\
transfusions of cryoprecipitate, platelets, fresh frozen plasma, and factor VII | 0\
chest was closed | 0\
severe cardiogenic shock | 24\
multiorgan failure | 24\
hypotensive | 24\
vasopressin | 24\
epinephrine | 24\
norepinephrine | 24\
hypoxic respiratory failure | 24\
mechanical ventilation | 24\
liver failure | 24\
albumin | 24\
blood products | 24\
broad-spectrum antibiotics | 24\
oliguric | 24\
continuous venovenous hemodialysis | 24\
acute renal failure | 24\
bilateral, symmetrical cyanotic changes to all 5 digits of his upper and lower extremities | 48\
vasopressor administration was stopped | 48\
surface pallor and coldness in the affected areas | 48\
upper- and lower-digit ischemia had progressed to dry gangrene | 216\
dull pain | 216\
no ability to move his fingers and toes | 216\
bilateral stiffness | 216\
2+ pitting edema | 216\
nonexistent capillary refill time | 216\
palpable 2+ peripheral pulses | 216\
Doppler study showed flat waveforms on all digits and toes bilaterally | 216\
no proximal occlusion or stenosis | 216\
intra-aortic balloon pump was removed | 168\
endotracheal tube was removed | 168\
albumin was discontinued | 264\
liver enzymes returned to normal limits | 264\
kidney function gradually improved | 984\
hemodialysis was stopped | 984\
mental status improved | 984\
necrotic lesions were treated conservatively with povidone-iodine dressings | 984\
debridement | 648\
negative-pressure wound therapy | 648\
purulent, foul-smelling material from his left infraclavicular operative site | 648\
stabilized and transferred to our facility | 1296\
laser extraction of his retained lead | 1392\
pus was drained from the subfascial area within the infraclavicular space | 1392\
antibiotic regimen | 1392\
microbial cultures grew Enterobacter cloacae and Staphylococcus epidermidis | 1392\
screening for subcutaneous implantable cardioverter-defibrillator | 1392\
transvenous implantable cardioverter-defibrillator system was implanted | 1536\
evaluation of his hands and feet revealed no signs of local infection or wet gangrene | 1536\
black skin changes and demarcation lines were clearly defined | 1536\
frank mummification of his digits and toes | 1536\
discharged to home health services | 1848\
amputation and debridement of his necrotic feet | 2544\
amputation of his fingers is scheduled | 2544