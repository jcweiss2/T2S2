six-year-old | 0
22.4kg | 0
female | 0
admitted to the pediatric intensive care unit | 0
febrile illness | -216
shortness of breath | -48
acute hypoxic respiratory failure | 0
septic shock | 0
suspected pneumonia | 0
diffuse bilateral interstitial opacities | 0
non-invasive positive pressure ventilation | 0
tracheal intubation | 6
empiric broad spectrum antibiotics | 0
sedation | 0
tidal volume 200ml | 0
respiratory rate of 30 | 0
PEEP of 6 cmH2O | 0
FiO2 1.0 | 0
mean airway pressure 21 cmH2O | 0
peak inspiratory pressure 32 cmH2O | 0
oxygenation index 19.3 | 0
PaO2:FiO2 ratio 102.3 | 0
severe PARDS | 0
arterial blood gas analysis | 0
pH 7.27 | 0
PaCO2 49 | 0
PaO2 87 | 0
base deficit 4.8 | 0
prone positioning | 0
paralysis | 0
worsening chest x-ray | 6
transthoracic echocardiogram | 6
normal function | 6
LV shortening fraction 54.9% | 6
no signs of pulmonary hypertension | 6
esophageal balloon catheter | 6
transpulmonary pressure measurement | 6
optimal titration of PEEP | 6
esophageal balloon placement | 6
gentle pressure applied to the abdomen | 6
cardiac oscillations detected | 6
thoracic ribcage pressure increase | 6
optimal positioning of the esophageal balloon | 6
PL ≤ 10 cm H2O | 6
PLexp 0 ± 2 cmH2O | 6
tidal volume titration | 6
PEEP titration | 6
neuromuscular blockade discontinued | 72
weaning PEEP | 72
esophageal balloon removed | 103
stable PLexp | 103
extubated | 155
weaned off respiratory support | 155