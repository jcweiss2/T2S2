29 years old | 0
Asian | 0
female | 0
gravida 1 | 0
para 0 | 0
admitted to the hospital | 0
fever | -216
nasal discharge | -216
coughing | -216
prescribed antibiotics | -216
admission due to orthopnoea | 0
exacerbation of respiratory distress | 0
wet-warm clinical phenotype of heart failure | 0
systolic murmur | 0
bilateral coarse crackles | 0
bilateral leg oedema | 0
history of hypothyreosis | 0
levothyroxine treatment | 0
no intravenous drug use | 0
no cardiovascular diseases | 0
no congenital heart disease | 0
no rheumatic fever | 0
no valvular heart disease | 0
no malignancy | 0
no autoimmune disease | 0
no coagulation abnormalities | 0
no gestational hypertension | 0
no diabetes | 0
sinus tachycardia | 0
complete right branch bundle block | 0
massive pulmonary congestion | 0
elevated brain natriuretic peptide | 0
elevated C-reactive protein | 0
elevated white blood cell count | 0
severe mitral valve regurgitation | 0
mobile vegetations on mitral leaflets | 0
severe pulmonary hypertension | 0
left ventricular ejection fraction 71% | 0
normal ultrasound and non-stress test for foetus | 0
infective endocarditis suspected | 0
simultaneous emergent caesarean section and mitral valve replacement | 0
intramuscular injection of betamethasone | -5
caesarean section | 0
male infant delivered | 0
APGAR scores 1, 5, and 6 | 0
uterine compression suture | 0
biological valve replacement | 0
mitral valve leaflets occupied by vegetations | 0
anterior mitral leaflet perforation | 0
histopathological examination of mitral valve | 24
acute neutrophil-dominant inflammation | 24
empiric intravenous antibiotic therapy | 0
extubation | 24
cardiac rehabilitation | 24
left ICU for general ward | 24
occlusion of mid-left anterior descending artery | 168
occlusion of peripheral right coronary artery | 168
multiple asymptomatic cerebral infarctions | 168
discharged | 696
neonate discharged | 4560
one-year follow-up echocardiography | 8760
normal mitral valve function | 8760
slightly decreased left ventricular ejection fraction | 8760