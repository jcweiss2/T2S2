59 years old | 0
female | 0
admitted to the hospital | 0
type-1 diabetes | -24000
end-stage renal failure | -24000
combined kidney-pancreas transplant | -24000
second kidney transplant | -8400
mycophenolate mofetil | -8400
tacrolimus | -8400
immunosuppressive regimen | -8400
10-day course of intravenous antibiotics | -240
no clinical improvement | -240
bilateral pleural effusion | 0
bilateral pneumonia | 0
multiple abdominal intussusceptions | 0
discontinued immunosuppressive treatment | 0
exploratory laparotomy | 0
free intra-abdominal liquid | 0
4 sites of intussusception | 0
intramural lesion | 0
post-transplant lymphoproliferative disorder | 0
biopsy of one of the lesions | 0
manual desinvagination | 0
low-grade tubulovillous adenoma | 0
new episode of bowel obstruction | 288
CT scan | 288
1 intussusception | 288
progression of pulmonary infection | 288
second surgery | 288
recurrence of the intussusception | 288
manual reduction of the invagination | 288
no clinical improvement | 288
multiple organ failure | 294
death | 294
autopsy | 294
multiple tubulovillous adenomas | 294
massive necrosis of the pancreas graft | 294
thrombosis of the pancreatic artery | 294
pulmonary adenocarcinoma | 294
multiple bilateral pulmonary metastases | 294
lymphangitic carcinomatosis | 294