62 years old | 0
male | 0
admitted to the hospital | 0
COVID-19 | -72
dyspnea | -72
asthenia | -72
cough | 0
fever | 0
oxygen saturation 93% | 0
hypertension | 0
left hydronephrosis | 0
kidney stones | 0
bilateral pneumonia | 0
diffuse ground-glass opacity | 0
nasal intermittent positive pressure ventilation | 0
Venturi mask | 0
oxygen at 14 l/m | 0
continuous positive airway pressure | 0
endotracheal intubation | 24
mechanical ventilation | 24
lung-protective ventilation | 24
prone position | 24
Klebsiella pneumoniae | 336
bronchoaspirate | 336
consolidation in the left lower lobe | 336
D-dimer increase | 336
Staphylococcus capitis | 504
Stenotrophomonas maltophilia | 504
bronchoaspiration | 504
severe hypoxemia | 504
ventilator maladjustment | 504
severe respiratory acidosis | 504
hypotension | 504
tracheostomy | 720
death | 888
postmortem lower respiratory tract swab for COVID-19 | 888
suppurative pericarditis | 888
mural thrombi | 888
superficial microhemorrhagic areas | 888
parenchymal congestion | 888
necrotic area | 888
liver parenchymal congestion | 888
glomerular collapse | 888
acute tubulointerstitial nephritis | 888
thrombosis of the renal arterioles | 888
hepatic centrilobular vein thrombosis | 888
periportal inflammation | 888
massive dilatation and congestion of the hepatic sinusoids | 888
mild cholestasis | 888
pulmonary fibrosis | 888
DAD | 888
vascular microthrombosis | 888
fibrosis with obliteration of the lumen | 888
parenchymal cells | 888
fibroblasts | 888
macrophages | 888
type II hyperplastic pneumocytes | 888