65 years old | 0
man | 0
diet-controlled type 2 diabetes mellitus | 0
hyperlipidemia | 0
stage 3 chronic kidney disease | 0
cardiac arrest | -17520
presented to the emergency department | -48
chills | -96
body aches | -96
shortness of breath | -96
cough productive of yellow sputum tinged with blood | -96
denied sick contacts | -96
denied travel in the past 2 years | -96
no hospitalizations in the preceding 6 months | -4320
heavy alcohol use | -17520
smoking prior to 2014 | -17520
confused | -48
hypoxemic | -48
chest radiograph consolidation right mid-lung | -48
azithromycin | -48
ceftriaxone | -48
did not improve on supplemental oxygen | -24
intubated | -24
blood cultures grew non-lactose fermenting Gram-negative rods | -24
respiratory cultures grew non-lactose fermenting Gram-negative rods | -24
meropenem | -24
levofloxacin | -24
amikacin | -24
lymphopenia | 0
persistent elevation in blood lactate | 0
worsening thrombocytopenia | 0
acute kidney injury | 0
high oxygen requirements despite mechanical ventilation | 0
repeat chest radiograph progression of disease | 0
transferred to ICU | 0
extracorporeal membrane oxygenation support | 0
septic shock unresponsive to 3 vasopressors | 0
chest auscultation coarse breath sounds | 0
lower extremities cool and mottled | 0
digits cool and mottled | 0
100% oxygen necessary to maintain saturations above 88% | 0
Acinetobacter baumannii identified in respiratory cultures | 0
Acinetobacter baumannii identified in blood cultures | 0
sensitive to all antimicrobials tested | 0
therapy narrowed to cefepime | 0
repeat cultures negative | 0
persistent lactic acidosis | 0
disseminated intravascular coagulopathy | 0
AKI necessitating hemodialysis | 0
bullae observed on legs | 240
dry gangrene on digits | 240
family requested withdrawal of life support | 264
expired | 264
