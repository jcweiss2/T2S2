62 years old | 0
    male | 0
    admitted to the hospital | 0
    brought to the emergency department | 0
    progressive shortness of breath | 0
    altered mental status | 0
    coronary artery disease | -35040
    drug-eluting stent implantation in the left anterior descending coronary artery | -35040
    hypertension | -35040
    hyperlipidemia | -35040
    diabetes mellitus | -35040
    chronic obstructive pulmonary disease | -35040
    alcoholism | -35040
    morbid obesity | -35040
    hypotensive | 0
    blood pressure 80/50 mm Hg | 0
    hypoxic respiratory failure | 0
    partial pressure of oxygen 76 mm Hg | 0
    emergently intubated | 0
    started on pressors | 0
    transferred to the intensive care unit | 0
    chest radiography bilateral infiltrates | 0
    right pleural effusion | 0
    electrocardiography normal sinus rhythm | 0
    new low voltage | 0
    old left-axis deviation | 0
    hyponatremia | 0
    acute kidney injury | 0
    leukocytosis | 0
    lymphopenia | 0
    mildly macrocytic anemia | 0
    coagulation panel within normal limits | 0
    elevated d-dimer | 0
    negative serial troponins | 0
    echocardiography large pericardial effusion | 0
    tamponade physiology | 0
    emergent pericardiocentesis | 0
    pericardial pressure 35 mm Hg | 0
    1.1 L of sanguinous fluid drained | 0
    right heart catheterization | 0
    sanguinous fluid | 0
    bloody sanguinous fluid | 0
    1.2 million red blood cells | 0
    cytology peripheral blood components only | 0
    no malignant cells | 0
    initial nasopharyngeal swab for COVID-19 negative | 0
    bronchoalveolar lavage sample positive for COVID-19 | 48
    drain output decreased | 120
    drain output stopped | 120
    repeat echocardiography resolution of pericardial effusion | 120
    drain removed | 120
    treated with hydroxychloroquine | 0
    treated with ribavirin | 0
    treated with lopinavir# 0.75x + 3 = 6, then x is

## Answers

Answered by

0

Answer:

x=4

Step-by-step explanation:

0.75x+3=6

0.75x=6-3

0.75x=3

x=3/0.75

x=4

Answered by

0

Answer:

x = 4

Step-by-step explanation:

0.75x + 3 = 6

0.75x = 6 - 3

0.75x = 3

x = 3 / 0.75

x = 4

hope it helps

please mark brainliest

Similar questions