32 years old | 0 | 0 
female | 0 | 0 
admitted to the hospital | 0 | 0 
fever | -168 | 0 
chills | -168 | 0 
generalized weakness | -168 | 0 
shortness of breath | -72 | 0 
intravenous drug use | -10080 | 0 
attention deficit/hyperactivity disorder | -10080 | 0 
dextroamphetamine/amphetamine | -10080 | 0 
abusing fentanyl intravenously | -10080 | 0 
non-smoker | 0 | 0 
does not consume alcohol | 0 | 0 
Temperature 102.7 °Fahrenheit | 0 | 0 
blood pressure 102/56 mmHg | 0 | 0 
pulse 136 beats per minute | 0 | 0 
respiratory rate 38 breaths per minute | 0 | 0 
oxygen saturation 94% on room air | 0 | 0 
moderate respiratory distress | 0 | 0 
bilateral rhonchi | 0 | 0 
tachycardia | 0 | 0 
no murmur, rub or gallop | 0 | 0 
white blood cell count (WBC) of 12,200/mm3 | 0 | 0 
hemoglobin of 10.9 g/dL | 0 | 0 
platelet count of 85,000/mm3 | 0 | 0 
ESR of 60 mm/hr | 0 | 0 
hyponatremia with a sodium of 124 mmol/L | 0 | 0 
creatinine level of 2.8 mg/dL | 0 | 0 
BUN of 98 mg/dL | 0 | 0 
NT-proBNP of 1028 pg/mL | 0 | 0 
sinus tachycardia | 0 | 0 
bilateral lower lobe infiltrates | 0 | 0 
small pleural effusions | 0 | 0 
given IV fluids | 0 | 24 
given levofloxacin intravenously | 0 | 24 
transferred to the intensive care unit | 24 | 24 
septic shock | 24 | 24 
acute respiratory failure | 24 | 24 
pressor support | 24 | 168 
mechanical ventilation | 24 | 168 
blood cultures grew gram-positive cocci | 24 | 24 
started on vancomycin therapy | 24 | 168 
large vegetation at the tip of anterior leaflet of tricuspid valve | 48 | 48 
moderate-to-severe tricuspid regurgitation | 48 | 48 
patent foramen ovale with shunt | 48 | 48 
multiple cavitary peripheral lung nodules | 48 | 48 
septic emboli | 48 | 48 
non-oliguric AKI | 48 | 168 
required renal replacement therapy | 48 | 168 
acute tubular necrosis | 48 | 168 
perfusion-related kidney injury | 48 | 168 
septic shock | 48 | 168 
MSSA | 72 | 72 
started oxacillin treatment | 72 | 168 
improved on supportive and antimicrobial therapy | 72 | 240 
weaned off pressors | 168 | 168 
successfully extubated | 168 | 168 
renal function started to recover | 168 | 240 
bilateral nontender purpuric papules | 240 | 240 
skin examination | 240 | 240 
bullous lesions | 264 | 264 
no mucosal or palmar involvement | 240 | 240 
no abdominal pain | 240 | 240 
no arthralgias | 240 | 240 
no paresthesia | 240 | 240 
no fever | 240 | 240 
no chills | 240 | 240 
HIV antibody negative | 240 | 240 
hepatitis B serology negative | 240 | 240 
p-ANCA negative | 240 | 240 
c-ANCA negative | 240 | 240 
cryoglobulin negative | 240 | 240 
rheumatoid factor negative | 240 | 240 
ANA weakly positive | 240 | 240 
anti-ds DNA antibody negative | 240 | 240 
Complement C3 low | 240 | 240 
Complement C4 normal | 240 | 240 
anti−HCV antibody positive | 240 | 240 
HCV viral load of 4.16 × 105 IU/mL | 240 | 240 
eosinophil count normal | 240 | 240 
aspirated fluid from her bullous lesions did not grow bacteria | 264 | 264 
no organisms seen on gram staining | 264 | 264 
punch biopsies from the bullous skin lesions showed perivascular neutrophil infiltration | 264 | 264 
fibrinoid necrosis of small vessels | 264 | 264 
leukocytoclastic vasculitis | 264 | 264 
no bacteria, fungi or evidence of viral inclusions | 264 | 264 
vancomycin started in lieu of oxacillin | 264 | 264 
progressive resolution of skin lesions | 264 | 312 
tricuspid valve replacement surgery | 312 | 312 
no perioperative complications | 312 | 312 
no recurrence of skin lesions | 744 | 744 
discharged | 744 | 744