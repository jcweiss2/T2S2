49 years old | 0
male | 0
presented to the emergency department | 0
one-week history of progressively worsening swollen scrotum | -168
one-week history of progressively worsening painful scrotum | -168
one-week history of progressively worsening swollen penis | -168
one-week history of progressively worsening painful penis | -168
diagnosed with infective episode of balanitis | -720
discharged with course of Ciprofloxacin | -720
pyrexial | 0
temperature of 39°C | 0
swollen tender scrotum | 0
swollen tender penis | 0
significant scrotal oedema | 0
no gangrenous patches | 0
no skin breaks | 0
raised white blood cell count of 25.1×109/L | 0
C-reactive protein of 269mg/L | 0
unremarkable urine dipstick | 0
blood cultures taken | 0
empirical antibiotics commenced | 0
intravenous Gentamicin | 0
intravenous Co-amoxiclav | 0
scrotal ultrasound scan revealed scrotal cellulitis | 0
scrotal ultrasound scan revealed oedema | 0
scrotal ultrasound scan revealed lymphadenopathy in the right inguinal canal | 0
CT thorax, abdomen, and pelvis performed | 0
no intra-abdominal pathology | 0
echocardiogram performed | 0
bilateral lower limb doppler study performed | 0
excluded infective endocarditis | 0
excluded deep vein thrombosis | 0
blood cultures revealed Streptococcus Anginosus | 0
antibiotics rationalised to Benzylpenicillin | 0
antibiotics rationalised to Clindamycin | 0
repeat ultrasound scan 3 days later | 72
demonstrated skin cellulitis | 72
suggested abscess in the root of the penis | 72
suggested abscess in the inguinal canal | 72
reactive hydroceles bilaterally | 72
concern regarding urethral involvement | 72
concern regarding ischiorectal involvement | 72
MRI performed same day | 72
MRI displayed 10×6cm abscess abutting ventral aspect of root of penis | 72
abscess extending to perineum | 72
abscess extending to base of scrotum | 72
displacing urethra | 72
not invading urethra | 72
incision and drainage of abscess undertaken in theatre | 72
returned to theatre for wound exploration and washout two days later | 168
third surgical exploration four days after initial surgery | 264
showed necrotic corpus cavernosum | 264
possible ischiorectal involvement | 264
flexible sigmoidoscopy showed normal recto-sigmoid colon up to 15cm | 264
suprapubic catheter sited | 264
comprehensive debridement of necrotic areas within corpora | 264
eight operative attempts at debridement | 264
eight operative attempts at wound washouts | 264
patient showed signs of clinical improvement | 264
antibiotic therapy continued for 5 weeks | 0
discharged after 6 weeks | 1008
declined to attend follow up | 1008
no information regarding reconstructive options | 1008
echocardiogram performed |1
bilateral lower limb doppler study performed |1
excluded infective endocarditis |1
excluded deep vein thrombosis |1
excluded infective endocarditis |
