male | 0
24 years old | 0
admitted to the hospital | 0
bilateral lumbago | -336
fever | -336
hematuria | -336
reduced urine volume | -336
gross hematuria | -336
visited another hospital | -336
no significant pain relief | -336
highest body temperature | 0
37.7 °C | 0
white blood cell | 0
42.08 × 10^9/L | 0
neutrophil count | 0
0.89 | 0
C-reactive protein | 0
271.42 mg/L | 0
procalcitonin | 0
46.97 ng/mL | 0
creatinine | 0
199 μmol/L | 0
Na | 0
123 mmol/L | 0
alanine aminotransferase | 0
63 U/L | 0
aspartate transaminase | 0
96 U/L | 0
total bilirubin | 0
177.3 μmol/L | 0
abscess drainage culture | 0
positive | 0
blood culture | 0
negative | 0
MRSA | 0
sensitive to vancomycin | 0
MIC 0.5 μg/mL | 0
vancomycin treatment | 0
1 g every 12 h | 0
CT scan | 0
multiple lesions | 0
inflammation | 0
abscess formation | 0
pneumatosis | 0
multiple calculi | 0
left kidney | 0
calculus | 0
left upper ureter | 0
mild dilation | 0
effusion | 0
left renal pelvis | 0
callyx | 0
upper ureter | 0
transferred to ICU | 120
fever | 120
shortness of breath | 120
respiratory rate | 120
33 bpm | 120
stable circulation | 120
fast heart rate | 120
116 bpm | 120
imipenem | 120
1 g every 8 h | 120
cilastatin sodium | 120
1 g every 8 h | 120
pathogenic metagenomics testing | 144
Streptomyces aureus | 144
presence | 144
blood | 144
right gluteus maximus drainage fluid | 144
culture | 144
MRSA | 144
sensitive to vancomycin | 144
MIC 1.5 μg/mL | 144
persistent hyperpyrexia | 168
highest temperature | 168
38.9 °C | 168
duration | 168
13 h | 168
new abscess | 168
anterior side | 168
left leg | 168
red | 168
swollen | 168
flowing liquid | 168
B-ultrasonography | 168
CT scans | 168
new infectious lesions | 168
decreases in inflammation indicators | 168
not significant | 168
CRP | 168
139.62 mg/L | 168
WBC | 168
26.86 × 10^9/L | 168
NEUT % | 168
0.883 | 168
daptomycin | 168
0.5 g daily | 168
linezolid | 168
0.6 g every 12 h | 168
treatment | 168
lung infection | 168
possible MRSA infection | 168
ultrasound-guided catheter drainage | 168
left renal pelvis | 168
fever | 192
persisted | 192
peak temperature | 192
38.8 °C | 192
duration | 192
10 h | 192
infection indicators | 192
lower | 192
CRP | 192
79.86 mg/L | 192
WBC | 192
19.17 × 10^9/L | 192
NEUT % | 192
0.841 | 192
PCT | 192
0.61 ng/mL | 192
stable respiration | 312
circulation | 312
shorter fever duration | 312
8 h | 312
decreased levels | 312
infection indicators | 312
transferred back | 312
general ward | 312
combination treatment | 312
daptomycin | 312
linezolid | 312
imipenem | 312
cilastatin sodium | 312
de-escalated | 312
cefoperazone sodium | 312
sulbactam sodium | 312
gram-negative bacteria infection | 312
culture | 432
negative | 432
no fever | 432
PCT | 504
0.21 ng/mL | 504
WBC | 504
10.36 × 10^9/L | 504
CRP | 504
35.56 mg/L | 504
NEUT % | 504
0.706 | 504
no fever | 504
stable condition | 504
discharged | 504
left nephrostomy tube | 504
unobstructed | 504
treated | 504
after complete recovery | 504