68 years old | 0
female | 0
hypothyroidism | 0
bipolar disorder | 0
sodium valproate | -7200
clozapine | -7200
risperidone | -7200
trihexyphenidyl | -7200
drowsy | -24
limb weakness | -24
hypothermic | -24
pulse 50/min | -24
blood pressure 90/60 mmHg | -24
respiratory rates 24/min | -24
bilateral plantars mute | -24
crepitations over right lower lung fields | -24
pancytopenia | -24
normal renal function | -24
normal liver function | -24
right lower and middle lobe consolidation | -24
crystalloids | 0
antibiotics | 0
hydrocortisone | 0
sepsis | 0
right lower zone pneumonia | 0
thyroid functions done | 0
thyroid-stimulating hormone 22.86 mIU/L | 0
normal FT4 | 0
normal FT3 | 0
anti-thyroid peroxidase antibodies negative | 0
thyroxine dose escalated | 0
respiratory distress worsened | 72
drowsy | 72
intubated | 72
mechanical ventilation | 72
vasopressors | 72
sedatives tapered | 168
infection brought under control | 168
vasopressors stopped | 168
lethargic | 168
poor respiratory efforts | 168
percutaneous tracheostomy | 240
magnetic resonance imaging brain normal | 240
cerebrospinal fluid examination normal | 240
total creatine kinase levels normal | 240
electroencephalography normal | 240
fixed gaze | 240
limited blinking | 240
fixed flexor posturing | 240
increased muscle tone | 240
psychiatry opinion | 240
provisional diagnosis of catatonia | 240
lorazepam test | 240
rigidity improved | 240
intravenous lorazepam | 240
fully conscious | 336
weaned off ventilator | 576
tracheostomy tube removed | 576
stoma strapped | 576
discharged | 840
doing well | 4320