16 years old | 0
female | 0
45 kg in weight | 0
157 cm in height | 0
left maxillary fracture | 0
no history of pulmonary disease | 0
no special features in electrocardiography | 0
no special features in biochemical examination of blood | 0
no special features in chest X-ray | 0
midazolam injection | -1
vital signs before anesthesia | -1
blood pressure 110/66 mmHg | -1
heart rate 80 beats/min | -1
oxygen saturation 99% | -1
induction of anesthesia with propofol | 0
loss of consciousness | 0
injection of rocuronium | 0
positive pressure ventilation | 0
tracheal intubation | 0
insertion of Mallinckrodt tube | 0
no leakage in the tube cuff | 0
normal breathing sound | 0
tidal volume and respiration rate maintained | 0
peak inspiratory pressure | 0
no air leakage | 0
anesthesia maintained | 0
oral irrigation with povidone iodine | 0
bubbles formed | 0
additional air inserted into the cuff | 0
bubbles continued to form | 0
tube removed | 0
povidone iodine drawn through a suction catheter | 0
tracheal intubation retaken | 0
new Mallinckrodt tube inserted | 0
normal breathing sound from both lungs | 0
pulse oxygen saturation 100% | 0
lung compliance and chest movement normal | 0
oral irrigation resumed | 0
no air leakage | 0
maximum inspiratory pressure | 0
oxygen saturation declined | 0.5
rale heard from the right lung | 0.5
operation stopped | 0.5
tracheal suction commenced | 0.5
frothy discharge came out | 0.5
chest X-ray conducted | 0.5
invasive arterial catheter inserted | 0.5
arterial blood gas analysis | 0.5
salbutamol nebulized | 0.5
methylprednisolone and furosemide injected | 0.5
mechanical ventilation with PEEP | 0.5
aspiration pneumonia in the right lung | 0.5
arterial blood gas analysis | 1
improvement in the patient's condition | 1
operation resumed | 1
operation finished | 1.5
pyridostigmine and glycopyrrolate used | 1.5
reversal of muscle relaxation | 1.5
spontaneous respiration recovered | 1.5
brownish-tinged liquid discharged | 1.5
suction through the tube | 1.5
povidone iodine aspirated | 1.5
trachea and bronchi cleaned with sterile saline solution | 1.5
fiberoptic bronchoscopy | 1.5
compliance of the reservoir bag improved | 1.5
arterial blood gas analysis | 1.5
patient transferred to intensive care unit | 2
mechanical ventilation continued | 2
antibiotics administered | 2
steroids and diuretics used | 2
tidal volume insufficient | 2
mechanical ventilation at pressure support mode | 2
arterial blood gas analysis | 7
leukocyte counts increased | 7
neutrophils increased | 7
body temperature increased | 7
fever diagnosed | 7
augmentin and cefepime prescribed | 7
methylprednisolone and furosemide administered | 7
pressure support and PEEP readjusted | 7
arterial blood gas analysis | 20
weaning performed | 25
T-piece used | 25
oxygen provided | 25
blood pressure and heart rate normal | 25
oxygen saturation remained high | 25
consciousness clear | 25
removal of the tube | 27
arterial blood gas analysis | 27
oxygen provided through nasal cannula | 27
arterial blood gas analysis | 32
oxygen saturation remained high | 32
oral discharge decreased | 32
chest X-ray showed improvement | 50
patient transferred to general ward | 50