54 years old | 0
Hispanic | 0
female | 0
type 2 diabetes | -8760
hypertension | -8760
peripheral vascular disease | -8760
right-foot transmetatarsal amputation | -26280
lisinopril | -72
metoprolol succinate | -72
pravastatin | -72
aspirin | -72
hydrochlorothiazide | -72
metformin | -72
insulin detemir | -72
insulin lispro | -48
severe watery diarrhea | -72
nausea | -72
vomiting | -72
mental status change | -72
hypoglycemia | 0
glucose level of 47 mg/dL | 0
glucagon administration | 0
confusion | 0
hypotension | 0
blood pressure of 70/39 mmHg | 0
disorientation | 0
dry oral mucosa | 0
decreased bowel sounds | 0
cardiopulmonary arrest | 0
pulseless electrical activity | 0
cardiopulmonary resuscitation | 0
endotracheal intubation | 0
mechanical ventilation | 0
norepinephrine | 0
vasopressin | 0
profound acidemia | 0
arterial pH 6.57 | 0
HCO3- 2 mEq/L | 0
anion gap 30 mmol/L | 0
osmolar gap of 21 | 0
lactate 16.3 mmol/L | 0
glycosylated hemoglobin 7.3 mg/dL | 0
creatinine of 8.07 mg/dL | 0
computed tomography scan of the abdomen and pelvis | 0
non-specific gallbladder wall thickening | 0
sepsis | 0
septic shock | 0
acute coronary event | 0
cardiogenic shock | 0
metformin toxicity | 0
renal replacement therapy | 0
hemodialysis | 0
continuous veno-venous hemofiltration | 0
type IV respiratory failure | 0
shock | 0
acidemia | 0
metformin concentration | 168
discontinuation of norepinephrine | 96
discontinuation of vasopressin | 96
extubation | 144
discharge from the intensive care unit | 216
discharge from the hospital | 360
gastroenteritis | -168
nuclear stress test | 360
coronary angiography | 360
three-vessel disease | 360
90% stenosis in the mid-left anterior descending artery | 360
80% stenosis in the first obtuse marginal artery | 360
90% stenosis in the mid-right coronary artery | 360
coronary artery bypass graft | 360
decreased level of consciousness | 0
lactic acidosis | 0
metformin-associated lactic acidosis | 0
acute kidney injury | 0
severe metabolic acidosis | 0
renal failure | 0
dialysis | 0
metformin use | -72
hypovolemia | 0
acute kidney injury | 0
gastrointestinal symptoms | 0
nausea | -72
vomiting | -72
abdominal pain | 0
leukocytosis | 0
mesenteric ischemia | 0
sepsis | 0
shock | 0
failure of standard supportive measures | 0
extracorporeal treatment | 0
lactate > 20 mmol/L | 0
pH 7.0 | 0
decreased level of consciousness | 0
metformin concentration | 168
troponin leak | 0
demand ischemia | 0
stable coronary artery disease | 0
profound metabolic and post-resuscitative hemodynamic stress | 0
elevated troponin of 4.42 ng/mL | 0
serial electrocardiograms | 0
echocardiogram | 48
ejection fraction of 50% | 48
regional wall motion abnormalities | 48
dialysis discontinuation | 720
renal function return to baseline | 720