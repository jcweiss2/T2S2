52 year old woman | 0
    high risk AML | -720
    recurrent Clostridioides difficile infection | -720
    admitted for one month prior | -720
    match-unrelated donor hematopoietic stem cell transplant | -720
    reduced intensity fludarabine-melphalan | -720
    tacrolimus | -720
    methotrexate | -720
    sepsis | -720
    metabolic encephalopathy | -720
    chronic diarrhea | -720
    transaminitis | -720
    acute kidney injury | -720
    bone graft failure | -720
    seen by infectious diseases in consultation several times | -720
    febrile neutropenia | -720
    encephalopathy | -720
    Klebsiella bacteremia | -720
    J. hoylei bacteremia | -720
    afebrile | 0
    normotensive | 0
    blood pressure 143/104 | 0
    pulse 104 beats per minute | 0
    respiratory rate 22 breaths per minute | 0
    oxygen saturation 97% | 0
    diffuse anasarca | 0
    bruising throughout extremities | 0
    bleeding gums | 0
    oral ulcers | 0
    mucositis | 0
    course bilateral breath sounds | 0
    hypoactive bowel sounds | 0
    oral mucosa without thrush | 0
    left chest PICC site clean | 0
    thirty days post-transplant | 0
    one aerobic blood culture | 0
    J. hoylei grew after 2 days and 20 hours | 0
    peripheral line | 0
    episode of decompensation | 0
    active oral mucositis hemorrhage | 0
    transferred to intensive care unit | 0
    airway management | 0
    organism grew on sheep blood agar after 48 hours | 0
    aerobic incubation at 37°C | 0
    5% CO2 | 0
    Gram-positive | 0
    coryneform | 0
    MALDI-TOF MS identification | 0
    16S ribosomal RNA gene PCR/sequencing | 0
    intravenous cefepime | -192
    vancomycin | -264
    empirically transitioned to imipenem | 0
    linezolid | 0
    ceftriaxone MIC >2 µg/mL | 0
    meropenem MIC ≤0.25 µg/mL | 0
    penicillin MIC 2 µg/mL | 0
    vancomycin MIC ≤1 µg/mL |%234