54 years old | 0
male | 0
admitted to the hospital | 0
motor vehicle collision | -1
Glasgow Coma Scale 13 | 0
intubated | 0
admitted to the surgical intensive care unit | 0
C1 transverse foramen fracture | 0
bilateral rib fractures | 0
pulmonary contusions | 0
febrile | 8
lower respiratory culture consistent with polymicrobial pneumonia | 48
started on broad-spectrum antibiotics | 48
significant active crack cocaine use | -24
quetiapine 400 mg at bedtime | -672
mirtazapine 30 mg at bedtime | -672
persistent intermittent agitation | 24
opioids | 24
dexmedetomidine | 24
lorazepam | 24
intravenous haloperidol 5 mg | 120
fever 102.2°F–104.7°F | 144
tachycardia | 144
hypertension | 144
diffuse lead-pipe rigidity | 144
hyperreflexia | 144
two-beat clonus | 144
differential diagnosis broadened to include sepsis, NMS, serotonin syndrome, and cocaine withdrawal | 144
serum creatine kinase 247 IU/L | 144
IV dantrolene 2.5 mg/kg | 144
quetiapine discontinued | 144
mirtazapine discontinued | 144
haloperidol discontinued | 144
dysautonomia resolved | 144.5
rigidity resolved | 144.5
hyperreflexia resolved | 144.5
temperature downtrended | 144.5
maintenance oral dantrolene | 168
resolution of rigidity | 168
improvement in fever curve | 168
bromocriptine added | 192
dantrolene discontinued | 360
rigidity recurred | 384
hyperreflexia recurred | 384
dantrolene restarted | 384
tapered 14-day course | 384
spontaneous breathing trial passed | 432
extubated | 432
mental status returned to baseline | 528
no further recurrence of symptoms | 528
quetiapine 50 mg QHS resumed | 528
discharged | 696