54 years old | 0
male | 0
admitted to the hospital | 0
ventral hernia | -720
increased in size | -168
became stony, hard, painful, and irreducible | -168
vomiting | -168
absolute constipation | -168
road-traffic accident | -7200
dysarthria | -7200
socially inactive | -7200
dehydrated | 0
pulse rate of 104 beats/minute | 0
blood pressure within normal range | 0
huge ventral hernia | 0
skin discoloration | 0
bowel sounds not audible | 0
rectal examination unremarkable | 0
leukocytosis | 0
chest x-ray showed no air under the diaphragm | 0
abdominal x-ray showed dilated bowel loops with few air fluid levels | 0
diagnosis of strangulated ventral hernia | 0
resuscitated with isotonic fluids | 0
intravenous cefuroxime and metronidazole | 0
operation | 2
laparotomy | 2
constriction at the abdominal wall | 2
pressure over the mesentery | 2
hernial sac opened | 2
offensive fluid and gangrenous bowel, mesentery, and omentum | 2
gangrenous area included most of the jejunum, as well as the entire ileum, cecum, and the ascending and proximal half of the transverse colon | 2
constriction divided | 2
trial to regain viability of the gut | 2
viability of the gut not regained | 2
decision to resect the gangrenous bowel and omentum | 2
resection of gangrenous bowel and omentum | 2
only 60 cm of proximal jejunum remained | 2
primary anastomosis | 2
direct hernia repair without prosthetic mesh | 2
histopathology showed gangrenous bowel with clear margins | 2
postoperative course uneventful | 2
total parenteral nutrition (TPN) started | 2
gradually overlapped with enteral feeding | 2
episodes of diarrhea managed conservatively | 2
discharged from the hospital | 720
short bowel syndrome | 720
followed in the outpatient surgical clinic | 720
combination of enteral and normal diet | 720
passing mixed-consistency stool 4 to 5 times a day | 720
lost approximately 30 kg of weight | 720
dietary issues managed with the help of a dietitian | 720