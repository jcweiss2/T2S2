54 years old | 0
female | 0
admitted with acute abdomen | 0
possible diagnosis intestinal obstruction | 0
required central line insertion | 0
central line insertion attempted under USG guidance in right subclavian vein | 0
started complaining of irritation near right ear | 0
guidewire inserted | 0
right IJV visualized under USG | 0
hyperechoic object seen | 0
guidewire confirmed in IJV | 0
guidewire taken out till not visible in IJV | 0
reattempts done while keeping probe over right IJV | 0
using routine methods putting pressure supraclavicular | 0
moving head toward right side | 0
assuring position of J point toward right atrium | 0
catheter inserted over guidewire | 0
guidewire removed | 0
venous aspiration from all three ports done | 0
saline flushed through catheter | 0
immediate turbulence in right atrium observed using microconvex probe | 0
catheter tip position in superior vena cava confirmed | 0
