89 years old | 0
male | 0
Caucasian | 0
admitted to the hospital | 0
fever | -168
cough | -168
warfarin | -4320
bisoprolol | -4320
ramipril | -4320
furosemide | -4320
valvular heart disease | -4320
atrial fibrillation | -4320
hypertension | -4320
SARS-CoV-2 infection | -240
amoxicillin | -240
spiramycin | -216
azithromycin | -192
epistaxis | 0
major bleeding | 0
hypoxaemia | 0
systolic blood pressure 105 mmHg | 0
diastolic blood pressure 59 mmHg | 0
cardiac rate 104 per minute | 0
INR > 10 | 0
D-dimers 400 ng/mL | 0
B-type natriuretic peptide 81 pg/mL | 0
high-sensitivity troponin T 10 ng/L | 0
ground-glass opacity | 0
crazy paving | 0
air space consolidation | 0
vitamin K 10 mg | 0
simple compression therapy | 0
liver injury ruled out | 0
fibrinogen level 7.6 g/L | 0
plasma D-dimer level 400 ng/mL | 0
antithrombin activity normal | 72
protein C chromogenic activity normal | 72
free protein S antigen normal | 72
G20210A F2 variant absent | 72
G1691A F5 variant absent | 72
antiphospholipid antibodies negative | 72
dexamethasone 6 mg per day | 0
cefotaxime | 0
azithromycin | 0
oxygen therapy | 0
INR fluctuations | 72
vitamin K administrations | 72
enoxaparin 100 IU/kg | 144
D-dimer increase > 12 000 ng/mL | 168
pulmonary embolism | 168
CTPA | 168
NT-proBNP 2022 ng/L | 168
high-sensitivity troponin T 48.9 ng/L | 168
tinzaparin 175 IU/kg | 216
discharged from ICU | 432
nasal oxygen therapy 2 L/min | 432
bacterial pneumonia | 480
septic shock | 576
death | 576
low-molecular-weight heparin therapy | 432
CYP2C9*2 variant | -4320
-1639G>A VKORC1 variant | -4320