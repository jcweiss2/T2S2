31 years old | 0
male | 0
admitted to the hospital | 0
severe abdominal pain | 0
tachycardia | 0
analgesics | 0
ERCP | 0
small rupture at the point where the fistulous tract joined the abdominal wall | 0
contrast material leaking into the abdominal cavity | 0
endoscopic sphincterotomy | 0
biliary stent placement | 0
fever | 48
diaphoresis | 48
tachycardia | 48
leucocytosis | 48
acute abdomen | 48
severe generalized biliary-purulent peritonitis | 48
hemodynamic instability | 48
bacteremia | 48
severe respiratory distress | 48
systemic inflammatory response syndrome | 48
septic shock | 48
multiresistant Pseudomonas aeruginosa | 48
discharged | 672
laparoscopic cholecystectomy | -672
CBD exploration | -672
T-tube placement | -672
uneventful postoperative course | -672
follow-up visit | -672
cholangiogram | -672
no contraindications for removal of the T-tube | -672
removal of the T-tube | -672
abdominal ultrasound | 0
small fluid collection | 0
conservative management | 24
ERCP | 24
abdominal lavage | 48
placement of abdominal drains | 48
sutured rupture of the fistulous tract | 48
intensive care unit admission | 48
ventilatory support | 48
multiple antibiotics | 48
vasoactive agents | 48
activated C protein | 48
