79 years old | 0
female | 0
abdominal pain | -672
nausea | -672
weight loss | -672
postprandial abdominal pain | -288
femoral–tibial bypass | -288
constipation | -288
discharged | -288
abdominal symptoms | -168
hemodynamic compromise | -168
distal superior mesenteric artery occlusion | -168
mucosal wall changes | -168
acute bowel ischemia | -168
peripheral vascular disease | 0
coronary artery disease | 0
asthma | 0
rheumatoid arthritis | 0
hypertension | 0
hyperlipidemia | 0
type 2 diabetes | 0
hypothyroidism | 0
breast cancer | 0
smoking history | 0
septic shock | 0
abdominal peritonitis | 0
hypoxemia | 0
hypotension | 0
anterior territory ST-segment elevations | 0
elevated troponin level | 0
SMA embolectomy | 0
resuscitation | 0
SMA thromboembolectomy | 0
resection of necrotic jejunum | 0
thromboembolic material | 0
pathologic examination | 0
intraoperative transesophageal echocardiography | 0
thrombus in pulmonary veins | 0
thrombus in left atrium | 0
biventricular dysfunction | 0
vasopressor support | 0
cardiac catheterization | 24
stenosis of right coronary artery | 24
stenosis of great saphenous vein bypass graft | 24
abdominal surgeries | 24
bowel resection | 24
spindle cell carcinoma of lung | 24
chest imaging | 24
mass in right upper lobe | 24
intraluminal thrombus burden | 24
pulmonary veins | 24
left atrium | 24
palliative measures | 336
diagnosis of spindle cell carcinoma | 168
postoperative complications | 168