46 years old | 0
    male | 0
    admitted to the hospital | 0
    left hip periprosthetic infection | 0
    sepsis | -24
    increased pain in the left hip | -24
    drainage of blood | -24
    purulence | -24
    open wound | -24
    no history of trauma in the left hip | 0
    no preceding fevers | 0
    no chills | 0
    severe psoriatic arthritis | 0
    steroids treatment | -672
    methotrexate treatment | -72
    left metal-on-metal THA | -157248
    right metal-on-metal THA | -78768
    elevated white blood cell count | 0
    decreased hemoglobin | 0
    decreased hematocrit |$|