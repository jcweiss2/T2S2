71 years old | 0
female | 0
admitted to the hospital | 0
acute loss of consciousness | 0
hypoglycemia | 0
swelling of left hand | 0
heat of left hand | 0
redness of left hand | 0
bite wound at tip of left middle finger | 0
dementia | -672
intravenous cefazolin | 0
cellulitis | 0
infection progression despite antibiotic treatment | 48
MRSA | 48
Kanavel’s cardinal signs of flexor tenosynovitis | 48
vancomycin infusion | 48
wound debridement | 48
partial amputation at distal interphalangeal joint | 48
decompression of median nerve | 48
purulent abscess | 48
redness persisted | 48
swelling persisted | 48
infection progression reduced | 48
abdominal pain | 120
dark brown blood in stool | 120
gastrointestinal bleed | 120
systemic shock | 120
systolic blood pressure 60 mmHg | 120
vasopressors administration | 120
elevated WBC count | 120
increased CRP | 120
increased creatinine | 120
reduced sodium | 120
reduced blood glucose | 120
reduced hemoglobin | 120
non-occlusive mesenteric ischemia | 120
emergency small bowel resection | 120
tube feedings | 120
norepinephrine addition | 120
SARS-CoV-2 exposure | 168
positive nasal swab test for COVID-19 | 168
acute pneumonia | 192
lung consolidation | 192
bilateral pleural effusions | 192
favipiravir treatment | 192
transfer to ICU | 192
hypervolemia | 192
increased oxygen demand | 192
continuous hemodiafiltration | 192
necrotizing fasciitis | 192
septic shock | 192
mechanical respiration | 192
high flow oxygen administration | 192
remdesivir treatment | 192
hydrocortisone administration | 192
osteomyelitis | 216
Vancomycin for osteomyelitis | 216
ARDS | 216
DIC | 240
ART-123 administration | 240
necrosis of entire third digit | 240
skin necrosis | 240
fascia necrosis | 240
musculature necrosis up to radio-carpal joint | 240
infection progression to forearm | 240
COVID-19 recovery | 336
mechanical ventilation weaning | 336
endotracheal tube withdrawal | 336
negative SARS-CoV-2 antigen test | 336
major amputation at distal third of forearm | 336
tissue debridement | 336
lavage | 336
heavy calcification of arteries | 336
tortuosity of arteries | 336
possible occlusions | 336
distal hypoperfusion ischemic syndrome | 336
skin flap coverage achieved | 336
stump closure | 336
septic shock recurrence | 672
cardiopulmonary arrest | 672
death | 672
