66 years old | 0
female | 0
endometrial cancer | 0
chemotherapy with doxorubicin and cisplatin | -192
neutropenic fever | 0
pancytopenia | 0
admitted to the hospital | 0
treated with broad-spectrum antibiotics | 0
hypoxic respiratory failure | 72
intubation | 72
endotracheal tube diameter, 8.0 mm | 72
acute pulmonary edema | 72
septic shock | 72
minute ventilation suddenly dropped | 72
mildly blood-tinged material | 72
suctioning the endotracheal tube | 72
chest radiography showed no change | 72
chest radiography showed a completely opacified left hemithorax | 84
no breath sounds over the left chest | 84
platelets were 38,000/µL | 84
flexible bronchoscopy | 84
large blood clot obstructing the proximal left main bronchus | 84
bronchoscopic lavage | 84
forceps extraction | 84
bronchoscopic cryotherapy | 84
blood clot frozen for 10 seconds | 84
blood clot removed in four large pieces | 84.25
follow-up chest X-ray | 84.25
significant improvement in aeration of the left lung | 84.25
no further obstructive events | 84.25
repeat bronchoscopic evaluation | 360
no evidence of the clot | 360
all of the airways were patent | 360
recovered from septic shock | 576
discharged from hospital | 576