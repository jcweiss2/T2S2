male | 0
preterm infant | 0
born at 28 weeks of gestation | 0
birth weight 1240g | 0
respiratory distress syndrome | 0
nasal continuous positive airway pressure | 0
caffeine citrate for apnoea of prematurity | 0
preterm formula started | 0
expressed breast milk | 0
feedings advanced | 0
increased gastric residual | -168
apnoea | -168
grossly bloody stools | -168
abdominal distention | -168
left abdominal tenderness | -168
sluggish bowel sounds | -168
increased C-reactive protein | -168
decreased white blood cell | -168
positive stool occult blood | -168
pneumatosis intestinalis | -168
feeds stopped | -168
intravenous antibiotics started | -168
pale and less active | -144
episodes of tachycardia and hypotension | -144
conventional mechanical ventilation | -144
fluid resuscitation | -144
haemodynamic support | -144
NEC diagnosis | -144
blood culture positive for Escherichia coli | -120
vancomycin stopped | -120
antibiotics changed | -120
conventional mechanical ventilation continued | -120
clinical and radiological improvement | -96
feedings resumed with expressed breast milk | -96
second episode of bloody stools | -24
abdomen soft | -24
non-tender | -24
active bowel sounds | -24
stool test positive for occult blood | -24
normal CRP and WBC levels | -24
mild thickening of the small bowel | -24
no evidence of pneumatosis intestinalis | -24
antibiotic therapy started | -24
feeding suspended | -24
serial blood analysis showed normal CRP and WBC levels | -18
enteral feeding with breast milk resumed | -18
antibiotics suspended | -18
third episode of bloody stool | 0
feeding with expressed mother’s milk fortified with cow’s milk | 0
infant quite well | 0
no emesis or abdominal distension | 0
active bowel sounds | 0
decreased WBC levels | 0
normal CRP levels | 0
mild increase in eosinophil counts | 0
FPIES suspected | 0
feeding suspended | 0
symptoms disappeared | 0
expressed mother’s milk fortified without cow’s milk | 0
no bloody stools | 0
preterm formula feeding reinitiated | 8
abdominal distension | 8
reoccurrence of grossly bloody stools | 8
normal WBC and CRP levels | 8
eosinophil count increased | 8
FPIES suspected | 8
formula changed to hydrolyzed formula | 8
resolution of symptoms | 8
discharged home | 60
breastfed for 8 months | 720
no recurrence of bloody stools | 720