14 years old | 0
African-American | 0
male | 0
admitted to the hospital | 0
right thigh pain | -24
painful ambulation | -24
no fever | -24
healthy | -24
no significant past medical history | -24
no trauma | -24
pain upon doing butterfly stretches | -24
mild leukocytosis | -24
erythrocyte sedimentation rate (ESR) of 10 mm/h | -24
C-reactive protein (CRP) of 5.7 mg/dL | -24
computed tomography (CT) of his pelvis | -24
magnetic resonance imaging (MRI) of the pelvis | -24
intramuscular tears | -24
edema | -24
mild widening of the right pubic bone apophysis | -24
osteitis pubis | -24
discharged | -24
crutches | -24
600 mg ibuprofen | -24
avoid sports | -24
follow-up with sports medicine | -24
readmitted to the hospital | 96
worsening symptoms | 96
abdominal pain | 96
thigh pain | 96
inability to walk | 96
worsening pain in both shoulders | 96
generalized myalgias | 96
malaise | 96
emesis | 96
diarrhea | 96
tachycardia | 96
tachypnea | 96
afebrile | 96
normotensive | 96
limited range of motion at the right hip | 96
diffuse tenderness to palpation | 96
no focal neurologic deficits | 96
white blood cell count of 12,100/µL | 96
ESR of 59 mm/h | 96
CRP of 20.7 | 96
CT of the abdomen and pelvis | 96
right obturator internus muscle fluid collection | 96
empirically given 1 gram of ceftriaxone | 96
started on intravenous vancomycin | 96
admitted to the intensive care unit | 96
oxacillin | 96
clindamycin | 96
blood and urine cultures | 96
urine cultures showed no growth | 96
blood cultures yielded methicillin sensitive Staphylococcus Aureus (MSSA) | 120
vancomycin discontinued | 120
MRI of the left shoulder | 120
repeat MRI of the pelvis | 120
myositis in the left shoulder | 120
enlarging fluid mass in the right obturator internus muscle | 120
osteomyelitis of the right pubic bone | 120
abscess drainage | 168
peripherally inserted central catheter (PICC) | 168
IV antibiotics | 168
Ancef 2 grams every 8 hours | 168
discharged | 216
denied any pain during ambulation | 216
white blood cells and ESR were noted to be 8900/µL and 79 mm/h | 216
physical therapy (PT) | 216
limitation in range of motion (ROM) | 224
strength from pain | 224
pressure present bilaterally at the anterior hips | 224
physical therapy proceeded | 224
gradual but significant improvement | 224
ESR and CRP gradually normalized | 224
peripherally inserted central catheter removed | 336
denied any pain with ambulation and climbing stairs | 336
full range of motion (ROM) and strength | 336
no further follow-up was needed | 336