6 years old | 0
female | 0
presented to the hospital | 0
right wrist swelling | -48
right wrist pain | -48
someone stepped on her wrist | -48
moderate pain | -48
worsened pain | -24
redness of the joint | -24
swelling of the joint | -24
subjective fever | -24
febrile | 0
tachycardic | 0
heart rate of 140 bpm | 0
swollen wrist | 0
erythematous wrist | 0
tender to palpation | 0
exquisite pain | 0
limited range of motion | 0
elevated ESR | 0
elevated CRP | 0
blood cultures drawn | 0
joint aspiration | 0
frankly purulent fluid | 0
gram-positive cocci | 0
numerous neutrophils | 0
IV clindamycin started | 0
admitted to the hospital | 0
arthrotomy | 24
seropurulent fluid | 24
joint space irrigated | 24
IV clindamycin continued | 24
afebrile | 48
pain well controlled | 48
repeat ESR | 48
repeat CRP | 48
joint aspiration fluid culture positive for Streptococcus pyogenes | 48
blood culture positive for Streptococcus pyogenes | 72
antibiotic regimen switched to IV cefazolin | 72
repeat arthrotomy | 96
no return of fluid | 96
joint irrigated and closed | 96
IV cefazolin continued | 96
serial ESR and CRP trended downward | 120
repeat blood culture showed no growth | 120
discharged | 144
oral cephalexin started | 144
ESR normalized | 240
CRP normalized | 240
completion of oral antibiotic course | 240