8.75 years old | 0
male | 0
neutered Burmese cat | 0
weighing 5.6 kg | 0
referred for treatment of pyothorax | 0
lethargy | -72
anorexia | -72
tachypnoea | -72
restrictive breathing pattern | -72
pyrexia | -72
bright | 0
alert | 0
responsive | 0
respiratory rate 40 breaths/min | 0
mild increase in respiratory effort | 0
heart rate 170 beats/min | 0
grade II/VI systolic murmur | 0
rectal temperature 38.1ºC | 0
hematocrit 36.3% | 0
WBCs 20.42 ×109/l | 0
neutrophils 17.97 ×109/l | 0
platelet count 185 ×109/l | 0
blood film analysis: mild neutrophilia with marked toxicity | 0
sodium 147 mmol/l | 0
potassium 4.1 mmol/l | 0
chloride 115 mmol/l | 0
calcium 1.31 mmol/l | 0
albumin 26 g/l | 0
globulin 34.6 g/l | 0
alanine aminotransferase 36.3 U/l | 0
total bilirubin 2.5 µmol/l | 0
creatinine 251 µmol/l | 0
urea 19 mmol/l | 0
creatinine kinase 1555 U/l | 0
lipaemia index none | 0
pH 7.292 | 0
PvCO2 44.2 mmHg | 0
glucose 8.9 mmol/l | 0
lactate 1.5 mmol/l | 0
HCO3– 19 mmol/l | 0
base excess -4.7 mmol/l | 0
USG 1.035 | 0
urine pH 6 | 0
urine protein 2+ | 0
urine culture negative | 0
pleural effusion analysis: neutrophilic septic exudate with intracellular cocci | 0
culture: beta-haemolytic Streptococcus agalactiae | 0
POCUS demonstrated pleural effusion | 0
thoracocentesis performed | 0
sedated with midazolam | 0
butorphanol | 0
alfaxalone | 0
bilateral chest drains placed | 0
thoracic radiographs taken | 0
thoracic drainage and lavage every 4h | 0
intrapleural bupivacaine 0.25% 1 mg/kg every 6h | 0
IV amoxicillin-clavulanate | 0
buprenorphine | 0
IV fluid therapy | 0
potassium chloride supplementation | 0
respiratory effort remained elevated 12h post-admission | 12
oxygen therapy initiated | 19
improvement in respiratory rate and effort 2h after initiating oxygen therapy | 21
FIO2 reduced to 0.4 | 21
oxygen therapy discontinued when respiratory parameters normalized | 19
mydriasis | 36
hypersalivation | 36
tonic-clonic seizure activity | 36
loss of consciousness | 36
sinus bradycardia 120 bpm | 36
blood pressure decreased to 110 mmHg systolic | 36
acidaemia pH 7.125 | 36
PvCO2 62.8 mmHg | 36
hypokalaemia 3.5 mmol/l | 36
hyperglycaemia 11.6 mmol/l | 36
hyperlactataemia 4.8 mmol/l | 36
creatinine 180 µmol/l | 36
suspected bupivacaine overdose | 36
confirmed dose 10 mg/kg | 36
ILE 20% bolus initiated | 36.25
mentation improved | 36.25
ILE CRI initiated | 36.25
thoracic lavage with NaCl 0.9% | 36.25
HR 140 bpm | 36.5
BP 130 mmHg systolic | 36.5
HR 160 bpm | 37.17
resolution of hypersalivation | 37.17
resolution of mydriasis | 37.17
intrapleural bupivacaine discontinued | 36.25
thoracic lavage continued | 36.25
resolving acidaemia pH 7.330 | 39
PvCO2 44.5 mmHg | 39
hypokalaemia 3.4 mmol/l | 39
azotaemia 162 µmol/l | 39
hyperglycaemia 8.3 mmol/l | 39
hyperlactataemia resolved | 39
mental status decline | 46
bradycardia 120-130 bpm | 46
second ILE bolus and CRI administered | 46.17
improved mentation | 46.17
bradycardia unresolved | 46.17
normotensive 140 mmHg systolic | 46.17
gradual improvement in mentation and HR | 56
oxygen therapy weaned over 44h | 80
general anaesthesia and CT performed | 76
right middle lung lobe abscess identified | 76
median sternotomy performed | 76
multiple episodes of hypotension | 76
treated with noradrenaline CRI | 76
respiratory distress secondary to laryngeal oedema | 76
re-intubated | 76
dexmedetomidine CRI initiated | 76
dexmedetomidine CRI discontinued | 79
analgesia tapered | 79
respiratory parameters normalized | 80
discharged on day 6 | 144
