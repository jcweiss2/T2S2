39 years old | 0
male | 0
documentary director | 0
living independently at home with his wife | 0
presented to the emergency department | 0
complaining of one-week long progressive epigastric pain | -168
associated nausea | -168
vomiting | -168
constipation | -168
past medical history of rectal adenocarcinoma | -9360
abdomino-perineal resection (APR) | -9360
end colostomy surgery | -9360
adjuvant chemoradiation therapy | -9360
non-smoker | 0
non-drinker | 0
septic shock | 0
fever | 0
temperature 39 °C | 0
tachycardic | 0
hypotensive | 0
BP 90/50 mmHg | 0
generalized abdominal tenderness | 0
guarding | 0
rebound tenderness | 0
leukocytosis | 0
anemia | 0
hemoglobin 8.6 mg/dL | 0
plain erect chest X-ray showed free air in the peritoneum | 0
nil by mouth | 0
septic management pathway activated | 0
IV fluid resuscitation | 0
IV broad-spectrum antibiotics | 0
pneumoperitoneum | 0
preliminary diagnosis of generalized peritonitis | 0
emergency laparotomy | 0
ileum perforated | 0
purulent fluid in the peritoneal cavity | 0
surgically resected | 0
anastomosis performed | 0
abdominal cavity wash out | 0
transferred to the intensive care unit | 0
close observation and monitoring | 0
hemodynamically unstable | 0
broad antibiotics (Imipenem, Tazocin, Vancomycin) | 0
antifungal medication (Caspofungin) | 0
continuous norepinephrine infusion | 0
fentanyl for pain and sedation | 0
continuous maintenance IV fluid therapy | 0
cardiac arrest | 36
resuscitated with CPR | 36
intensive fluid resuscitation | 36
extubated on day 5 post-op | 120
deteriorating clinically | 168
febrile | 168
triple (IV, oral, enema) contrasted abdominal CT | 168
large collection in the spleen containing gas and oral contrast | 168
colo-splenic fistula | 168
splenectomy | 168
left hemicolectomy | 168
moderately differentiated adenocarcinoma in splenic flexure of the colon | 168
extensive necrosis with foci of viable adenocarcinoma in the spleen | 168
uneventful recovery | 208
return of intestinal peristalsis | 208
increase in appetite | 208
resolved septic status | 208
discharged 40 days post-op | 960
followed up regularly at one-month | 1080
three-month | 1440
six-month | 2160
surveillance colonoscopy | 8760
ulcerated mass in the right colon | 8760
biopsy confirming adenocarcinoma | 8760
total colectomy and end ileostomy insertion | 8760