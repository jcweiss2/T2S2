30 years old | 0
woman | 0
bilateral liposuction | -10
unbearable pain in bilateral thigh liposuction sites | -10
erythema | -10
blisters | -10
admitted to our hospital | 0
febrile (38.2°C) | 0
heart rate of 128 beats/minute | 0
small scattered incisions in bilateral waist and thigh regions | 0
local skin over bilateral thighs exhibited swelling | 0
local skin over bilateral thighs exhibited tenderness | 0
blisters in posterior thigh region | 0
sutures removed in bilateral thigh regions |2 0
urine was black | 0
leukocytosis (25 ×10^9 cells/L) | 0
elevated C-reactive protein level (35 mg/dL) | 0
elevated serum creatinine level (250 U/L) | 0
elevated blood urea nitrogen level | 0
fasciotomy | 0
drainage of bilateral thighs | 0
treated with vancomycin | 0
treated with meropenem | 0
vital signs unstable | 0
diagnosed with sepsis | 0
diagnosed with renal insufficiency | 0
diagnosed with shock | 0
transferred to surgical intensive care unit | 0
continuous renal replacement therapy | 0
anti-infection treatment | 0
blood transfusion | 0
shock correction | 0
large amount of exudation in both thighs | 24
local swelling in both thighs | 24
extensive fasciotomy | 24
osteofascial compartment incision | 24
vacuum sealing drainage (VSD) of bilateral thigh regions | 24
degeneration of subcutaneous fat | 24
necrosis of subcutaneous fat | 24
degeneration of fascia | 24
necrosis of fascia | 24
degeneration of muscle | 24
necrosis of muscle | 24
