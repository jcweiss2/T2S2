71 years old | 0
male | 0
admitted to the hospital | 0
atrial fibrillation | -24
hospital admission for atrial fibrillation catheter ablation | -24
ostium secundum atrial septal defect | -24
mitral regurgitation | -24
atrial fibrillation catheter ablation | -24
transcatheter ostium secundum atrial septal defect repair | -24
discharged | -18
hospital admission for atrial fibrillation recurrence | 0
left atrial mass | 0
anticoagulant optimization | 0
apixaban to acenocoumarol | 0
persistent left atrial mass | 4
surgical removal of the mass | 4
left atrial myxoma | 4
last follow-up | 12
clinically stable | 12
permanent atrial fibrillation | 12
good echocardiographic surgical result | 12
no tumour recurrence | 12
pulmonary vein ablation | -24
transoesophageal echocardiography | -24
osASD | -24
significant left-to-right shunt | -24
coronary angiography | -24
no significant disease | -24
discharged on apixaban | -18
external electrical cardioversion | 0
physical examination unremarkable | 0
completely asymptomatic | 0
tranthoracic echocardiography | 0
moderate mitral regurgitation | 0
device-related thrombus | 0
acenocoumarol | 0
optimal intensity of anticoagulation | 0
TEE | 4
size of the mass unchanged | 4
isoechoic aspect | 4
irregular margins | 4
extreme mobility | 4
severe mitral regurgitation | 4
cardiovascular magnetic resonance imaging | 4
T1 isointensity | 4
T1 fat-saturated isointensity | 4
T2 hyperintensity | 4
first-pass perfusion enhancement absent | 4
late contrast enhancement difficult to assess | 4
coronary angiography | 4
neovascularization | 4
multidisciplinary heart team discussion | 4
cardiac surgery indicated | 4
LA mass resection | 4
closure device removal | 4
LA septum reconstruction | 4
pericardial patch | 4
mitral valve replacement | 4
bioprosthesis | 4
bileaflet prolapse | 4
macroscopic examination | 4
gelatinous surface | 4
friable surface | 4
irregular edges | 4
histopathological diagnosis | 4
myxoma | 4
intensive care unit | 4
pneumonia | 4
septic shock | 4
acute kidney injury | 4
inpatient rehabilitation facility | 42
asymptomatic | 12
permanent AF | 12
good surgical result | 12
no tumour recurrence | 12