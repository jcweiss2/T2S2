39 years old | 0
    African American man | 0
    admitted to the hospital | 0
    HIV | -672
    HAART noncompliance | -672
    MSM | -672
    anal receptive intercourse | -672
    facial swelling | -336
    lip swelling | -336
    painful rash | -336
    facial rash | -336
    scalp rash | -336
    torso rash | -336
    perianal rash | -336
    bowel movement pain | -336
    bright red blood per rectum | -336
    denial of recent travel | 0
    denial of contact with sick persons | 0
    afebrile | 0
    warm to the touch | 0
    vesiculopustular patches | 0
    facial ulceration | 0
    scalp ulceration | 0
    anal coalescing lesion | 0
    anal crusting | 0
    purulent discharge | 0
    rectal exam refusal | 0
    normal electrolytes | 0
    normal blood urea nitrogen | 0
    normal creatinine | 0
    anemia | 0
    low leukocytes | 0
    normal neutrophils | 0
    normal lymphocytes | 0
    normal eosinophils | 0
    normal monocytes | 0
    normal basophils | 0
    low CD4 count | 0
    normal liver function | 0
    MPX DNA PCR positive | 0
    high HIV viral load | 0
    negative chlamydia | 0
    negative gonorrhea | 0
    negative HSV IgM | 0
    rectal thickening | 0
    rectal lumen obliteration | 0
    pericolonic mesenteric stranding | 0
    perianal fistulas | 0
    MPX infection | 0
    proctitis | 0
    tecovirimat | 0
    Biktarvy | 0
    MPX vaccine declined | 0
    PEG | 0
    parenteral opiates | 0
    tramadol | 0
    gabapentin | 0
    blood transfusion | 0
    Bactrim | 0
    Azithromycin | 0
    deterioration | 24
    facial swelling persisted | 24
    rectal pain persisted | 24
    rash spreading | 24
    fever | 24
    Salmonella infection | 24
    Covid19 infection | 24
    MRSA infection | 24
    intravenous TPOXX | 24
    Vaccinia immunoglobulin | 24
    methylprednisolone | 24
    hypoxemic respiratory failure | 48
    ICU admission | 48
    bilateral pulmonary infiltrates | 48
    ARDS | 48
    septic shock | 48
    pneumonia | 48
    vasopressors | 48
    cardiac arrest | 48
    decreased cardiac function | 48
    sepsis | 48
    multiorgan failure | 48
    death | 48
    