48 years old | 0
male | 0
admitted to the hospital | 0
perianal abscess | 0
syphilis | -672
penicillin anaphylaxis | -672
routine blood tests | 0
Tolulized Red Unheated Serum Test | 0
etimiicin | -48
ornidazole | -48
incision and drainage | 0
neck pain | 1
dizziness | 1
chest pressure | 1
high blood pressure | 1
fever | 2
decreased blood pressure | 2
neutrophilic leukocytosis | 2
procalcitonin level | 2
fluid resuscitation | 2
temperature dropped | 2
transferred to ICU | 2
intravenous imipenem-cilastatin | 2
dopamine | 2
worsening neutrophilic leukocytosis | 48
procalcitonin value | 48
MODS | 72
abscess culture | 72
Neisseria gonorrhoeae | 72
Staphylococcus haemolyticus | 72
blood cultures | 72
R. mannitolilytica | 72
antibiotic therapy | 72
ceftriaxone | 72
levofloxacin | 72
repeat blood cultures | 144
no bacterial growth | 144
incision wound healed | 144
satisfactory recovery | 432
R. mannitolilytica infection | 0
sepsis | 2
multiple organ dysfunction syndromes | 72
bacteremia | 72
antimicrobial susceptibility | 72
minimum inhibitory concentration | 72
 MALDI-TOF Mass Spectrometry | 72
Bruker | 72
confidence level | 72
VITEK-2 CIMPACT | 72
broth microdilution method | 72
CLSI | 72
non-Enterobacteriaceae | 72
piperacillin/tazobactam | 72
cotrimoxazole | 72
quinolones | 72
third and fourth generation cephalosporins | 72
postoperative sepsis | 2
aminoglycosides | 2
Escherichia coli | 2
anuria | 2
elevated inflammatory markers | 2
dopamine | 2
broad-spectrum imipenem-cilastatin | 2
deep perianal infection | 2
pelvic magnetic resonance | 2
computed tomography | 2
abdomen | 2
chest | 2
multi-organ failure | 72
abnormal liver functions | 72
renal functions | 72
elevated cardiac enzymes | 72
bacterial culture | 72
drug sensitivity | 72
febrile patients | 72
opportunistic pathogens | 72
R. mannitolilytica infections | 0
immunocompromised patients | 0
immunocompromised person | 0
Treponema pallidum infections | 0
cellular immunity | 0
Th1/Th2 | 0
CD4+CD25− T cells | 0
CD4+ T cells | 0
CD4+/CD8+ | 0
gonorrhea | 72
sepsis | 2
opportunistic pathogen | 2
sensitive antibiotics | 72
culture results | 72
treatment guidelines | 72
drug susceptibility | 72
quinolones | 72
third and fourth generation cephalosporins | 72
piperacillin/tazobactam | 72
cotrimoxazole | 72
antibiotic therapy | 72
levofloxacin | 72
ceftriaxone | 72
S. haemolyticus | 72
N. gonorrhoeae | 72
syphilis spirochetes | 72
bacterial culture | 72
drug sensitivity | 72
febrile patients | 72
opportunistic pathogens | 72
R. mannitolilytica | 0
infections | 0
opportunistic pathogen | 0
multidrug-resistant profiles | 0
clinical practice | 0
treatment of infections | 0
opportunistic pathogens | 0
R. mannitolilytica | 0
 ethic approval | 0
consent to publish | 0
disclosure | 0