59 years old | 0
male | 0
hypertensive | 0
non-diabetic | 0
admitted to the hospital | 0
stapled hemorrhoidopexy | 0
rectal bleeding | -720
prolapsing piles | -720
metoprolol | -8760
amlodipine | -8760
4th degree piles | 0
large external component | 0
prophylactic antibiotics | -0.5
ceftriaxone | -0.5
gentamycin | -0.5
spinal anesthesia | 0
difficulty in closure | 0
hemorrhoids excised | 0
uneasiness | 0
discomfort | 0
midazolam | 0
hypotensive | 0
Ringer lactate | 0
tetrastarch | 0
stabilisation of mean arterial pressure | 0
fluid administered | 0
post-operative ward | 0
pain at the operative site | 2
butorphanol nasal spray | 2
generalized weakness | 24
breathlessness | 24
BP falling | 30
hypotension | 30
normal saline | 30
intensive care unit | 30.5
central line | 30.5
central venous pressure guided fluid therapy | 30.5
arterial blood gas analysis | 30.5
oxygen | 30.5
venturi mask | 30.5
non-invasive BP monitoring | 30.5
pulse rate monitoring | 30.5
heart rate monitoring | 30.5
SpO2 monitoring | 30.5
temperature monitoring | 30.5
continuous CVP monitoring | 30.5
urine output monitoring | 30.5
abdominal girth monitoring | 30.5
fever | 30.5
hypotension | 30.5
tachycardia | 30.5
respiratory distress | 30.5
decreased air entry | 30.5
fine crepts | 30.5
abdominal distension | 30.5
absent bowel sounds | 30.5
urinary catheterization | 30.5
sinus tachycardia | 30.5
noradrenaline | 30.5
dopamine | 30.5
metabolic acidosis | 30.5
low pO2 | 30.5
non-invasive biphasic positive airway pressure ventilation | 30.5
meropenem | 30.5
teicoplanin | 30.5
metronidazole | 30.5
urine output | 31
coagulation profile deranged | 31
fresh frozen plasma | 31
chest physiotherapy | 31
nebulization | 31
general nursing care | 31
hemodynamic parameters improved | 35
urine output improved | 35
ABG improved | 35
noradrenaline tapered | 35
dopamine tapered | 35
oxygen inhalation | 35
Hudson mask | 35
discharged | 216
rectal perforation | -720
peritonitis | -720
sepsis | 30
septic shock | 30
multi-organ failure | 30
mortality | -720
laparotomy | -720
fecal diversion | -720
low anterior resection | -720
rectal tissue excised | 0
bacterial entry | 0
peri-rectal sepsis | 30
retroperitoneal sepsis | 30
incomplete rings | 0
doughnuts | 0
excised rectal tissue | 0
sepsis treatment | 30
non-invasive ventilation | 30
antibiotics | 30
supportive care | 30
nursing care | 30