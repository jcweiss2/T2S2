38 years old | 0
female | 0
fever | -48
fatigue | -48
arthralgia | -48
furuncle-like skin lesion | -48
admitted to the hospital | 0
generalized abdominal pain | 0
nausea | 0
vomiting | 0
general discomfort | 0
nasogastric tube placement | 0
dyspnea grade IV | 0
desaturation | 0
CT scan | 0
right perirenal abscess | 0
thickening of the left renal vein | 0
bilateral pulmonary septic impacts | 0
bilateral mild pleural effusion | 0
bilateral hypoventilation | 0
jaundice | 0
oligoanuria | 0
low platelet count | 0
urine and blood cultures | 0
empirical treatment with vancomycin | 0
tazobactam | 0
anticoagulation treatment with Low Molecular Weight Heparin | 0
warfarin | 0
mechanical respiratory assistance | 0
dialysis | 0
clindamycin antibiotic | 0
fever persisted | 0
multi-organ failure | 0
blood culture positive for resistant methicillin staphylococcus | 12
gram negative bacillus in alveolar fluid wash | 12
vancomycin, daptomycin, and meropenem | 12
bacteremia | 12
persistent fever | 12
mechanical respiratory assistance with inotropic drugs | 12
new thorax abdomen and pelvis tomography | 12
phleboectasia | 12
extension of the thrombus | 12
surgical exploration | 12
informed consent | 12
bilateral nephrectomy | 12
torpid evolution | 24
feverish records | 24
colistin | 24
antibiotic scheme (vanco-dapto-mero-colistin) | 24
broncho alveolar lavage | 24
Serratia + Kleb KPC | 24
culture of intra-surgical samples show: Yeast | 24
fluconazole | 24
antibiotic scheme (vanco-dapto-mero-colistin-fluco) | 24
improvement | 35
antibiotic scheme (vanco-colistin-fluco) | 35
left thoracentesis | 35
antibiotic scheme (Vanco + Fluco + Colistin + Mero + Metronidazole) | 38
episodes of intermittently altered hemodynamic status | 38
vancomicine | 41
all other antibiotic suspended | 41
blood cultures | 41
adrenal profile | 41
suprarenal insufficiency | 41
hydrocortisone | 41
improved general condition | 41
transferred to the intermediate care unit | 63
discharged from hospital | 73
mental health follow-up | 73
awaiting a new evaluation for kidney transplantation | 73
decolonization treatment | 73
body cleaning per seven days with chlorhexidine | 73
daily application of mupirocin in the nostrils | 73