26 years old | 0\
male | 0\
admitted to the hospital | 0\
new-onset headache | 0\
blurred vision | 0\
kidney transplant | -6048\
end-stage kidney disease | -9120\
immunosuppression | 0\
mycofenolate sodium | 0\
methylprednisolone | 0\
estimated glomerular filtration rate (eGFR) | 0\
proteinuria | 0\
chronic kidney transplant disease | 0\
status post vascular rejection | -6048\
chronic calcineurin-inhibitor toxicity | -6048\
several contrast-enhancing intracerebral lesions | 0\
perifocal edema | 0\
methylprednisolone therapy stopped | 0\
dexamethasone | 0\
brain edema | 0\
transmitted to the university department of Nephrology | 0\
transmitted to the department of Neurosurgery | 0\
brain biopsy | 0\
cerebral PTLD | 0\
diffuse large B-cell lymphoma | 0\
positive for Ebstein-Barr virus | 0\
initial chemotherapy regime | 0\
high-dose cytarabin | 0\
Rituximab | 0\
complete remission of PTLD | 168\
impairment of the transplant function | 168\
eGFR | 168\
cytomegalovirus (CMV) reactivated | 336\
pneumocystis jirovecii pneumonia | 336\
chemotherapy changed to Rituximab | 336\
antiviral and antibiotic therapy | 336\
mycofenolate sodium tapered | 336\
generalized seizure | 720\
recurrence of PTLD | 720\
cerebral MRI scan | 720\
HDMTX | 720\
Leukovorine | 720\
Rituximab | 720\
vigorous hydration | 720\
HFHD | 744\
dialysis procedures | 744\
MTX-level in serum | 744\
no acute kidney failure | 744\
nadir of leucocytes | 780\
CMV- and E.coli pneumonia | 936\
sepsis | 936\
acute kidney transplant failure | 936\
transmission to an intensive care unit | 936\
invasive ventilation | 936\
sepsis managed | 936\
follow up cerebral MRI scan | 1096\
small regredience of PTLD | 1096\
cerebral radiation | 1096\
no relevant response of the disease | 1096