66 years old| 0
male | 0
fever | -288
cough | -288
arthralgia | -288
influenza-like illness | -288
diagnosed with type-A influenza | -288
oseltamivir | -288
high fever continued | -288
dyspnea gradually progressed | -288
admitted to a nearby hospital | -168
chest CT showed bilateral multiple granular shadows | -168
chest CT showed patchy opacities | -168
MRSA detected in sputum culture | -168
treated with sulbactam/ampicillin | -168
treated with levofloxacin | -168
CRP reduced from 40.0 to 23.0 mg/dL | -168
bilateral consolidation on chest X-ray worsened | -168
transferred to our hospital | 0
conscious | 0
temperature 38.2 ºC | 0
blood pressure 149/79 mmHg | 0
heart rate 118 beats/minute | 0
respiratory rate 20 breaths/minute | 0
oxygen saturation 98% under 3 L/min oxygen | 0
faint coarse crackles in bilateral lungs | 0
no wounds observed | 0
leukocytosis with predominant neutrophils | 0
hypoalbuminemia | 0
CRP elevated 19.14 mg/dL | 0
procalcitonin 2.43 ng/mL | 0
sIL-2R elevated 2,475.0 U/mL | 0
rheumatoid factor normal | 0
antinuclear antibodies normal | 0
anticytoplasmic antibodies normal | 0
chest X-ray showed bilateral infiltration | 0
chest CT showed multiple cavities | 0
chest CT showed surrounding ground-grass opacities | 0
chest CT showed bilateral pleural effusion | 0
treated with sulbactam/ampicillin | 0
performed bronchoscopy | 48
suctioning of purulent sputum | 48
biopsy | 48
brushing cytology | 48
gram staining showed gram-positive cocci | 48
cytological examination showed neutrophils with phagocytosis | 48
histopathological examination showed necrosis | 48
inflammatory exudate | 48
fibrin deposition | 48
immature fibrosis | 48
pulmonary abscesses | 48
treated with vancomycin 1,000 mg/day | 96
vancomycin increased to 1,500 mg/day | 96
MRSA sensitive to trimethoprim/sulfamethoxazole | 96
MRSA sensitive to erythromycin | 96
MRSA sensitive to minocycline | 96
MRSA sensitive to clindamycin | 96
MRSA sensitive to vancomycin | 96
type IV SCCmec identified | 96
PVL gene identified | 96
diagnosed with necrotizing pneumonia due to CA-MRSA | 96
vancomycin reduced temperature | 96
vancomycin reduced white blood cell count | 96
vancomycin reduced CRP | 96
oxygenation resolved | 96
pulmonary opacities improved | 96
changed to linezolid due to drug-induced fever | 648
sputum negative for MRSA | 720
sputum negative for bacteria | 720
discharged | 984
chest CT showed disappearance of cavities | 4320
farmer | 0
current heavy smoker 96 pack-years | 0
never traveled abroad | 0
no recent contact with foreigners | 0
history of pneumonia | 0
history of acute renal failure | 0
no medical problems until 12 days before admission | -288
not vaccinated for influenza | 0
no vegetation in cardiac valves | 0
no deep vein thrombosis | 0
no septic embolism | 0
no invasive pulmonary aspergillosis | 0
no cryptogenic organizing pneumonia | 0
no granulomatosis with polyangiitis | 0
no pulmonary malignancies | 0
blood cultures negative | 0
bilateral multiple consolidations improved | 720
cavities improved | 720
anti-MRSA agents stopped | 984
complete improvement of general condition | 984
Aspergillus antigen positive | 0
β-D-glucan 13.4 pg/mL | 0
CEA 2.1 ng/mL | 0
CA19-9 2.9 U/mL | 0
influenza A negative | 0
influenza B negative | 0
Mycobacterium tuberculosis negative | 0
cryptococcus antigen negative | 0
Candida antigen negative | 0
rheumatoid factor 5 U/mL | 0
ANA <x40 | 0
