72 years old | 0
hispanic | 0
male | 0
admitted to the hospital | 0
pulmonary fibrosis | -672
oral steroids | -672
home oxygen therapy | -672
hypertension | -672
diabetes mellitus | -672
no prior smoking history | -672
progressive dyspnea | -168
cough | -168
productive of yellow sputum | -168
no hemoptysis | -168
fever | -168
night sweats | -168
six-pound weight loss | -168
scalp lesion | -336
pain | -336
no pruritus | -336
no discharge | -336
temperature of 96.8°F | 0
blood pressure of 153/87 | 0
heart rate of 82 | 0
respiratory rate of 22 | 0
oxygen saturation of 86% | 0
ulcerative lesion | 0
cervical lymphadenopathy | 0
fine bilateral diffuse crackles | 0
leukocytosis | 0
white blood count of 23,200 Cells/mcL | 0
hemoglobin of 12.3 g/dL | 0
platelets of 211,000/mcL | 0
blood urea nitrogen of 17 mg/dL | 0
creatinine of 0.8 mg/dL | 0
arterial blood gas | 0
pH of 7.44 | 0
PO2 of 51 | 0
PCO2 of 39 | 0
gradient of 50 mmHg | 0
bilateral interstitial infiltrates | 0
intravenous corticosteroids | 0
oxygen | 0
nebulized treatments | 0
severe pulmonary hypertension | 24
echocardiogram | 24
diffuse fibrotic changes | 24
multiple densities | 24
CT-guided biopsy | 48
poorly differentiated malignant neoplasm | 48
foci of necrosis | 48
immunohistochemical stains | 48
adenocarcinoma | 48
genotype testing | 48
EGFR mutation | 48
RAS mutation | 48
alk translocation | 48
excision of the right scalp lesion | 72
poorly differentiated malignant neoplasm | 72
immunohistochemical stains | 72
severe hypoxic respiratory failure | 120
intubation | 120
transfer to the intensive care unit | 120
septic shock | 120
healthcare associated pneumonia | 120
vasopressors | 120
intravenous antibiotics | 120
deteriorated | 336
expired | 336