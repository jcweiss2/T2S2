65 years old | 0
    female | 0
    admitted to the hospital | 0
    fever | 0
    chills | 0
    pain in left leg | 0
    parkinsonism | -17520
    diabetes mellitus | -17520
    levodopa / carbidopa | -17520
    rasagiline | -17520
    ropinirole | -17520
    trihexyphenidyl | -17520
    amantadine | -17520
    metformin | -17520
    glipizide | -17520
    cellulitis | 0
    intravenous clindamycin | 0
    intravenous benzylpenicillin | 0
    high-temperature spikes | 72
    tachycardia | 72
    tachypnea | 72
    hypotensive | 72
    encephalopathic | 72
    shifted to ICU | 72
    sepsis with multi-organ dysfunction syndrome | 72
    intravenous linezolid | 72
    intravenous piperacillin with tazobactam | 72
    hemodynamics improved | 72
    minimal inotropic supports | 72
    oral hypoglycemic agents stopped | 72
    insulin started | 72
    confused | 72
    drowsy | 72
    disoriented | 72
    altered sensorium | 72
    myoclonus | 72
    tremors | 72
    jerky movements | 72
    no neck stiffness | 72
    computed tomography of the brain | 72
    cerebrospinal fluid analysis | 72
    improving white blood cell counts | 72
    better glycemic control | 72
    sterile blood and pus cultures | 72
    high temperature | 96
    altered mental status | 96
    myoclonus | 96
    jerky movements | 96
    tremors | 96
    rasagiline continued | 96
    linezolid started | 96
    serotonin syndrome suspected | 96
    linezolid stopped | 120
    rasagiline stopped | 120
    temperature settled | 128
    heart rate normal | 144
    sensorium improved | 144
    tremors subsided | 144
    shifted out of ICU | 168
    started walking with support | 240
    discharged | 240
    anti-parkinsonism drugs continued | 240
    rasagiline restarted | 240
    regular follow-up with neurologist | 240
    stable | 240
    asymptomatic for serotonin syndrome | 240

    