40 years old | 0
male | 0
admitted to the hospital | 0
diabetic | -8760
COVID-19 | -360
hospitalized | -360
medication | -360
ventilator support | -360
discharge from the hospital | -336
unilateral swelling | -336
loosening of teeth | -336
mucormycosis | -336
surgical debridement | -336
amphotericin B drug therapy | -336
oroantral communication | -336
oronasal communication | -336
mastication difficulties | -336
nasal regurgitations | -336
absence of the left orbit | -336
total maxilla | -336
concave profile | -336
nasolabial fold | -336
corners of mouth drooped | -336
insufficient upper lip support | -336
full complement of teeth | -336
porcelain-fused ceramic full-veneer crown | -336
supraerupted malaligned anterior teeth | -336
normal tongue | -336
normal temporomandibular joint movement | -336
left total maxillectomy | -336
right subtotal maxillectomy | -336
left orbital decompression | -336
resection of the left zygomatic arch | -336
resection of the left zygomatic rim | -336
implant-supported removable prosthesis | 0
custom-made subperiosteal zygomatic implants | 0
titanium | 0
surgical procedure | 0
general anesthesia | 0
implant placement | 0
abutments | 0
open-tray impression copings | 15
impression | 15
inter arch records | 15
aluminum-coated wax | 15
titanium metal bar | 15
obturator | 15
acrylic resin material | 15
prosthesis insertion | 15
postinsertion instructions | 15
denture instructions | 15
oral hygiene instructions | 15
heat-cured acrylic resin | 15
metal mesh | 15
bilateral balance occlusion | 15
semianatomic teeth | 15
polyvinyl siloxane impression materials | 15
follow-up visit | 24
reline | 24
soft relining material | 24
follow-up visits | 39
occlusal refinements | 39
speech quality | 39
peripheral seal | 39
patient satisfaction | 90
satisfied with prosthesis | 90