70 years old | 0
male | 0
laparoscopic abdominoperineal resection (APR) | 0
adjuvant chemotherapy with oxaliplatin | 0
adjuvant chemotherapy with fluorouracil | 0
adjuvant chemotherapy with calcium folinate | 0
perineal hernia | -10920
reconstruction of the pelvic floor with Permacol™ mesh | -10920
transperineal approach | -10920
postoperative course uneventful | -10920
pelvic–abdominal CT scan | -7800
no locoregional recurrence | -7800
no reherniation | -7800
weight loss | -1560
thoracic–abdominal CT scan | -1560
multiple liver metastases | -1560
multiple lung metastases | -1560
chemotherapy with bevacizumab | -1560
chemotherapy with irinotecan | -1560
chemotherapy with calcium folinate | -1560
chemotherapy with fluorouracil | -1560
sepsis signs | 0
high temperature | 0
tachycardia | 0
hypotension | 0
pain in right buttock | 0
infection signs at area | 0
acute US examination | 0
abscess revealed | 0
US-guided drainage | 0
intensive unit admission | 0
intravenous fluids | 0
broad-spectrum antibiotics | 0
CT scan with contrast | 0
subcutaneous abscess cavity in perineum | 0
communication to small bowel | 0
laparotomy | 0
perineal fistula from distal ileum | 0
small bowel resection | 0
primary anastomosis | 0
postoperative complications | 24
severe fluid disturbances | 24
severe electrolyte disturbances | 24
intensive care unit stay | 24
pressors treatment | 24
parenteral nutrition | 24
perineal wound vacuum-assisted closure | 168
discharge to hospice | 672
