35 years old | 0
female | 0
pregnant | 0
admitted to the hospital | 0
fever | -240
cough | -240
dyspnoea | -120
aggravated dyspnoea | -120
cyanosis of the lip | 0
thick breathing sounds in both lungs | 0
dry and wet rales in the right lower lung | 0
tachycardia | 0
respiratory rate of 20 times/min | 0
COVID-19 infection | -240
S. aureus infection | -240
respiratory failure | 0
pregnancy with 34 + 4 wk | 0
G2P1 | 0
left occiput anterior | 0
elderly second parturient women | 0
maternal lower weight | 0
oligohydramnion | 0
premature live baby | 0
electrolyte disturbance | 0
hypoproteinaemia | 0
caesarean section | 24
oxyhemoglobin saturation improved | 24
discharged from the hospital | 264
chest CT showed multiple plaques | 0
miliary foci | 0
nodular foci with partial consolidation and cavities | 0
obstetric ultrasound showed a single viable foetus | 0
head presentation | 0
oligohydramnios | 0
cardiac ultrasound and lower extremity vascular ultrasound showed no significant abnormalities | 0
metagenomic next-generation sequencing (mNGS) | 24
S. aureus combined with novel coronavirus infection | 24
antibiotic therapy | 24
anticoagulant therapy | 24
treatments to relieve the cough and reduce the amount of sputum | 24
symptomatic treatment | 24
nasal tube oxygen | 48
chest CT showed multiple areas of inflammation in both lungs | 96
mildly enlarged mediastinal lymph nodes | 96
small amount of bilateral pleural effusion | 96
CRP was 38.54 mg/L | 96
WBC count was 8.25 × 10^9/L | 96
PCT was 0.129 ng/mL | 96
potassium was 4.04 mmol/L | 96
D-dimer was 2.44 mg/L | 96
TB-PCR was negative | 96
antibiotics were adjusted to sitafloxacin | 216
patient was discharged from the hospital | 264
chest CT showed that the multiple lung inflammation was absorbed slightly | 288
chest CT showed that the multiple lung inflammation was apparently absorbed | 336
S. aureus was resistant to both macrolide and lincosamide antibiotics | 24
inflammatory lesions of the patients’ lungs were gradually absorbed and improved | 216