57 years old | 0
female | 0
no significant medical history | 0
habitual use of alcohol | 0
habitual use of tobacco | 0
habitual use of diet supplements | 0
fever | -72
diarrhea | -72
ingestion of tetracycline | -72
fatigue | -72
admitted to a local general hospital | -72
elevated transaminase levels | -72
bicytopenia | -72
reduced prothrombin time activity | -72
hepatitis A virus-specific IgM antibodies negative | -72
hepatitis B surface antigen negative | -72
hepatitis C virus antibody negative | -72
viral capsid antigen negative | -72
cytomegalovirus antigenemia negative | -72
antimitochondrial antibody negative | -72
anti-smooth muscle antibody negative | -72
HTLV-1 antibody negative | -72
HIV antibody negative | -72
encephalopathy | -72
confusion | -72
slow movement | -72
bone marrow biopsy | -72
increased numbers of maturity histiocytes | -72
hemophagocytosis | -72
diagnosed with fulminant hepatitis | -72
diagnosed with hemophagocytic syndrome | -72
steroid pulse therapy | -72
continuous hemodiafiltration | -72
transferred to our hospital | 0
severe respiratory failure | 72
tracheal intubation | 72
mechanical ventilation | 72
computed tomography of the chest | 72
bronchial wall thickening | 72
bilateral diffuse infiltration shadow of lungs | 72
bronchoscopic findings | 72
pseudomembranous formation | 72
β-D-glucan level increased | 72
Aspergillus galactomannan antigen positive | 72
C-reactive protein increased | 72
procalcitonin increased | 72
blood gas test | 72
pH | 72
PaO2 | 72
PaCO2 | 72
HCO3- | 72
PaO2/FiO2 | 72
endobronchial biopsy | 72
active inflammation | 72
necrotic tissue | 72
filamentous fungal hyphae infiltration | 72
Aspergillus fumigatus isolated | 72
Burkholderia cepacia isolated | 72
diagnosed with pseudomembranous ITBA | 72
diagnosed with acute respiratory distress syndrome | 72
broad-spectrum antibiotics | 72
antifungal therapy | 72
voriconazole | 72
caspofungin | 72
β-D-glucan level decreased | 120
tracheobronchial pseudomembrane scarring | 120
septic shock | 120
Burkholderia cepacia | 120
acute respiratory distress syndrome | 120
died | 1368