79 years old | 0
    lady | 0
    presented with occipital headache | -48
    nausea | -48
    vomiting | -48
    past medical history of herpes zoster infection | 0
    hypertension | 0
    hyperlipidemia | 0
    labyrinthitis | 0
    Ramsay Hunt syndrome | 0
    previous hysterectomy | 0
    tonsillectomy | 0
    breast operations | 0
    cataract operations | 0
    ramipril | 0
    bisoprolol | 0
    atorvastatin | 0
    clopidogrel | 0
    aspirin | 0
    zolpidem | 0
    alfacalcidol | 0
    calcium | 0
    no drug allergies | 0
    hyponatremia at 126 mmol/L | 0
    increased GGT 198 mmol/L | 0
    bilirubin 19 mmol/L | 0
    normal bloods | 0
    clear urinalysis | 0
    CT brain was normal | 0
    chest radiograph showed mild pulmonary vascular congestion | 0
    no chest pain | 0
    no abdominal pain | 0
    provisional diagnosis of encephalitis | 0
    antibiotics started | 0
    lumbar puncture refused on admission | 0
    lumbar puncture done on Day 4 | 96
    herpes simplex virus 1 infection | 96
    acyclovir commenced | 96
    ultrasound on Day 13 | 312
    nonspecific abdominal pain | 312
    cholelithiasis | 312
    no cholecystitis | 312
    conservative treatment continued | 312
    pain localized to the right iliac fossa | 336
    CT abdomen pelvis showed ischemia | 336
    pneumatosis | 336
    laparotomy on Day 18 | 432
    bowel ischemia | 432
    retrocaecal perforation | 432
    terminal ileal band | 432
    internal herniation | 432
    gangrene | 432
    extended right hemicolectomy | 432
    maximum dose of inotropes | 432
    abdominal wall kept open | 432
    Bogota bag | 432
    re-look surgery in 24 hours | 432
    no progression of ischemia | 456
    stabilized patient | 456
    ileostomy formed | 456
    closure of abdomen | 456
    spent 18 days in intensive care unit | 432
    bowel ischemia not due to sepsis | 432
    bowel ischemia not due to hypovolemia | 432
    innocent adhesional band | 432
    potentially life-threatening clinical condition | 432
    arterial phase CT abdomen pelvis | 336
    acute bowel ischemia of terminal ileum | 336
    acute bowel ischemia of ascending colon | 336
    pneumatosis | 336
    suspected hypoperfusion | 432
    long intensive care unit stay | 432
    mechanical cause found on laparotomy | 432
    terminal ileal band precipitated internal herniation | 432
    compromise of bowel | 432
    gangrene | 432
    retrocaecal perforation | 432
    surgical revascularization | 432
    resection of affected bowel | 432
    extended right hemicolectomy | 432
    ileostomy | 456
    aggressive fluid resuscitation | 432
    careful choice of vasoactive drugs | 432
    high level of suspicion needed | 0
    early surgical intervention | 432