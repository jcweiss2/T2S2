79 years old | 0
    female | 0
    diagnosed with acute pancreatitis | 0
    high fever | 0
    involuntary weight loss | 0
    inadequate nutrient consumption | 0
    two episodes of vomiting | 0
    severe pain in upper right abdomen | 0
    comorbid diabetes | 0
    hypertension | 0
    history of atrial fibrillation | -26208
    history of cholestasis | -26208
    underweight status | 0
    identified as at risk for refeeding syndrome | 0
    sudden pain | 0
    intense pain | 0
    nausea | 0
    lack of appetite | 0
    received ciprofloxacin | 0
    received metronidazole | 0
    elevated C-reactive protein concentration | 0
    elevated erythrocyte sedimentation rate | 0
    elevated leukocyte count | 0
    signs of inflammation around pancreas on computed tomography | 0
    no alcohol consumption | 0
    no organ failure | 0
    diagnosed with steatosis | 0
    diagnosed with cholelithiasis | 0
    refeeding as principal cause of rapid deterioration | 0
    poor oral intake | 0
    weight loss | 0
    pancreatitis contributing to refeeding syndrome | 0
    uncomfortable | 0
    sweating | 0
    wheezing | 0
    accelerated breathing | 0
    full mental awareness | 0
    dehydrated | 0
    pulse rate 90 beats/minute | 0
    blood pressure 135/75 mmHg | 0
    body temperature 38.5°C | 0
    no thoracic pathologic findings | 0
    modest mitral murmur | 0
    local tenderness in right upper abdomen | 0
    no muscular defense | 0
    positive Murphy sign | 0
    positive Blumberg sign | 0
    gallbladder enlargement | 0
    gallbladder stones | 0
    common bile duct expansion | 0
    pancreatic inhomogeneous echostructure | 0
    bile calculi | 0
    lack of appetite | 0
    reduced dietary intake for more than 5 days | 0
    low potassium concentration | 0
    low phosphate concentration | 0
    low magnesium concentration | 0
    respiratory failure | 0
    cardiac failure | 0
    treated with intravenous antimicrobial therapy | 0
    treated with intravenous rehydration therapy | 0
    treated with 0.5% glucose | 0
    treated with spasmolytic drugs | 0
    nutritional assessment | 48
    maintained oral feeding | 48
    retrograde endoscopic cholangiopancreatography | 72
    enteral feeding through nasogastric tube | 96
    refused oral feeding | 96
    low-speed normocaloric enteral feeding | 96
    enteral preparation | 96
    enteral feeding interrupted | 96
    confusion | 96
    tachycardia | 96
    respiratory insufficiency | 96
    severe hypotension | 96
    treated with rapid fluid supplementation | 96
    oxygen supplementation | 96
    treated with dopamine | 96
    severe electrolyte alterations | 96
    severe vitamin deficiencies | 96
    hydric balance dysfunction | 96
    diagnosed with refeeding syndrome | 96
    enteral feeding suspended | 96
    scheduled parenteral feeding | 96
    parenteral feeding bag insertion | 96
    mild recovery | 120
    started oral feeding | 120
    calorie intake 10 kcal/kg | 120
    phosphorus supplementation | 120
    potassium supplementation | 120
    magnesium supplementation | 120
    sodium supplementation | 120
    increased calorie intake by 5 kcal/kg | 168
    thiamine supplementation | 168
    increased calorie intake by 20-30 kcal/kg | 192
    monitored liver function | 192
    monitored kidney function | 192
    supplemented fluids | 192
    supplemented electrolytes | 192
    further increased calorie intake | 312
    clinical improvement | 312
    decreased body temperature to 36.8°C | 312
    normalized laboratory parameters | 312
    electrocardiogram no ischemia | 312
    echocardiogram low ejection fraction | 312
    bilateral pleural effusion | 312
    resumed small oral intake | 336
    stabilized hemodynamic status | 336
    discontinued vasopressor therapy | 336
    electrolyte imbalance disappeared | 336
    