muscle and joint pain | -144
general weakness | -144
fever | -144
liver dysfunction | -144
systemic inflammation | -144
admission | 0
continuous sedation | 0
muscle relaxation | 0
intubation | 0
mechanical ventilation | 0
broad-spectrum empirical antimicrobial therapy | 0
methylprednisolone | 0
stress ulcer prophylaxis | 0
thromboprophylaxis | 0
prone position | 0
chest CT | 0
bedside focus ultrasound | 12
acute renal failure | 144
CRRT | 144
CytoSorb adsorber installation | 168
septic episode | 240
second CytoSorb therapy session | 240
ICU delirium | 240
antipsychotics | 240
percutaneous tracheostomy | 240
weaning off from ventilator | 336
transfer to general ward | 1152
transfer to rehabilitation clinic | 1200
discontinuation of norepinephrine | 192
discontinuation of norepinephrine after second therapy | 264
decrease in CRP levels | 168
decrease in leukocyte levels | 168
improvement in ventilation parameters | 168
improvement in lung function | 168
reduction in extravascular lung water | 168
stabilization of pulmonary capillary integrity | 168
reduction in inflammation markers | 168
gradual improvement in patient condition | 168