36 years old| 0
    female | 0
    pregnant at 16 weeks and 1 day | 0
    lower abdominal pain | -24
    flank pain | -24
    vaginal spotting | -24
    mild dysuria | -24
    urinary frequency | -24
    urgency | -24
    no fever | -24
    no chills | -24
    no sick contacts | -24
    arrived in the United States from Pakistan | -5760
    blood pressure 103/70 mmHg | 0
    heart rate 133 bpm | 0
    temperature 99.9°F | 0
    respiratory rate 16 per minute | 0
    oxygen saturation 99% | 0
    well appearing | 0
    tachycardia | 0
    suprapubic tenderness | 0
    no rebound | 0
    no guarding | 0
    pelvic examination with slight bleeding | 0
    no uterine tenderness | 0
    leukocytosis 16.1 K/μL | 0
    88% polymorphonuclear leukocytes | 0
    normal complete blood count | 0
    normal chemistry panels | 0
    normal urinalysis | 0
    live intrauterine pregnancy | 0
    gestational age 16 weeks and 0 days | 0
    fetal heart rate 182 bpm | 0
    normal MRI abdomen | 0
    no appendicitis | 0
    received normal saline | 0
    received morphine sulfate | 0
    received acetaminophen | 0
    heart rate improved to 100 bpm | 0
    discharged home | 0
    returned to ED | 24
    sudden onset vaginal bleeding | 24
    abdominal pain | 24
    heart rate 139 bpm | 24
    blood pressure 149/88 mmHg | 24
    respiratory rate 30 per minute | 24
    oxygen saturation 100% | 24
    actively delivering products of conception | 24
    received misoprostol | 24
    tympanic temperature 105°F | 24
    persistent tachycardia into the 140s | 24
    hemodynamically unstable | 24
    blood pressure 84/35 mmHg | 24
    central intravenous access obtained | 24
    given acetaminophen | 24
    given normal saline | 24
    given vancomycin | 24
    given piperacillin/tazobactam | 24
    working diagnosis sepsis of unknown etiology | 24
    venous pH 7.22 | 24
    anion gap 21 | 24
    lactate concentration 10.8 mmol/L | 24
    white blood cell count 14.9 K/μL | 24
    85% polymorphonuclear leukocytes | 24
    normal MRI | 24
    normal urinalysis | 24
    no colitis | 24
    no skin infection | 24
    no soft tissue infections | 24
    given norepinephrine | 24
    admitted to medical intensive care unit | 24
    received ampicillin | 24
    received gentamycin | 24
    received clindamycin | 24
    suspected chorioamnionitis | 24
    ultrasonogram suggestive retained products of conception | 24
    underwent dilatation and curettage | 24
    removal of tissue debris | 24
    discharged from hospital | 96
    blood cultures positive H influenzae | 24
    retroplacental hemorrhage | 24
    placental abruption | 24
    adjacent infarct | 24
    no acute chorioamnionitis | 24
    spontaneous abortion | 24
    
    