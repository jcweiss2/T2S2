56 years old | 0
male | 0
obese | 0
smoker | 0
occasional alcohol drinker | 0
admitted to the Hospital Emergency Department | 0
oppressive holocranial headache | -120
fever | -120
hearing loss | -120
vomiting | -120
dysthermic sensation | -120
onset of the disease | -120
preparation, handling, and intake of roast pork | -120
anxiolytic (diazepam) | -120
analgesics (metamizole, tramadol) | -120
antiemetic (metoclopramide) | -120
persistent headache | 0
diaphoresis | 0
signs of meningeal irritation | 0
progressive state of agitation | 0
cranial computed tomography scan | 0
lumbar puncture | 0
cerebrospinal fluid (CSF) with a cloudy-whitish appearance | 0
white blood cell count 18.7 x 103/µL | 0
hemoglobin 15.2 g/dL | 0
platelet count 115 x 103/µL | 0
glucose 141 mg/dL | 0
creatinine 0.8 mg/dL | 0
lactate 15.7 mg/dL | 0
C-reactive protein 7 mg/dL | 0
procalcitonin 0.45 ng/mL | 0
CSF cytochemical characteristics | 0
glucose <10 mg/dL | 0
total protein 950 mg/dL | 0
13,720 leukocytes/µL | 0
Gram-positive diplococci | 0
admitted to the Intensive Care Unit (ICU) | 0
dexamethasone | 0
broad-spectrum antimicrobial therapy | 0
ampicillin | 0
ceftriaxone | 0
vancomycin | 0
acyclovir | 0
alpha-hemolytic streptococci isolation | 24
S. suis identification | 24
antibiotic resistance profile | 24
antibiotic susceptibility to penicillin | 24
antibiotic susceptibility to cefotaxime | 24
antibiotic susceptibility to levofloxacin | 24
antibiotic susceptibility to vancomycin | 24
antimicrobial targeted treatment with cefotaxime | 24
ICU admission | 0
favorable clinical evolution | 144
referred to the Internal Medicine Service | 144
audiometry | 168
complementary tests | 168
hearing loss exacerbation | 168
tinnitus | 168
discharged | 672
amoxicillin / clavulanic acid | 672
follow-up with the specialists | 672