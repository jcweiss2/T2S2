3 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
fever | -168 | 0 | Factual
diarrhea | -168 | 0 | Factual
abdominal pain | -168 | 0 | Factual
severe dehydration | -168 | 0 | Factual
admitted to the hospital | 0 | 0 | Factual
tachypneic | 0 | 0 | Factual
rapid shallow breathing | 0 | 0 | Factual
hypotensive | 0 | 0 | Factual
purpuric eruption | 0 | 0 | Factual
no organomegaly | 0 | 0 | Negated
no lymphadenopathy | 0 | 0 | Negated
pancytopenia | 0 | 0 | Factual
absolute neutropenia | 0 | 0 | Factual
renal impairment | 0 | 0 | Factual
electrolyte imbalance | 0 | 0 | Factual
hyperuricemia | 0 | 0 | Factual
coagulopathy | 0 | 0 | Factual
disseminated intravascular coagulation | 0 | 0 | Factual
high inflammatory markers | 0 | 0 | Factual
gram-negative Bacilli Escherichia coli | 0 | 0 | Factual
intravenous fluid therapy | 0 | 168 | Factual
blood components transfusion | 0 | 168 | Factual
correction of electrolyte disturbance | 0 | 168 | Factual
antibiotic therapy | 0 | 168 | Factual
provisional diagnosis of acute infectious gastroenteritis | 0 | 0 | Factual
sepsis | 0 | 0 | Factual
severe dehydration | 0 | 0 | Factual
acute renal failure | 0 | 0 | Factual
disseminated intravascular coagulation | 0 | 0 | Factual
discharged | 168 | 168 | Factual
unexplained irritability | 504 | 504 | Factual
abnormal behavior | 504 | 504 | Factual
hallucinations | 504 | 504 | Factual
failure to recognize parents | 504 | 504 | Factual
cerebral venous sinus thrombosis | 504 | 504 | Factual
thrombosis in both the left sigmoid and the transverse sinuses | 504 | 504 | Factual
low molecular weight heparin | 504 | 720 | Factual
improved | 720 | 720 | Factual
discharged | 720 | 720 | Factual
follow-up appointment | 720 | 720 | Factual
readmitted | 1008 | 1008 | Factual
fever | 1008 | 1008 | Factual
pallor | 1008 | 1008 | Factual
abdominal enlargement | 1008 | 1008 | Factual
leukocytosis | 1008 | 1008 | Factual
anemia | 1008 | 1008 | Factual
thrombocytopenia | 1008 | 1008 | Factual
blast cells | 1008 | 1008 | Factual
hepatosplenomegaly | 1008 | 1008 | Factual
bone marrow examination | 1008 | 1008 | Factual
hypercellular bone marrow | 1008 | 1008 | Factual
blast cells | 1008 | 1008 | Factual
immunophenotyping | 1008 | 1008 | Factual
diagnosis of Common ALL | 1008 | 1008 | Factual
induction therapy | 1008 | 1344 | Factual
consolidation | 1344 | 1680 | Factual
thrombophilia mutations panel | 1344 | 1344 | Factual
positive factor XIII V34L | 1344 | 1344 | Factual
MTHFR A1298C homozygous mutations | 1344 | 1344 | Factual
heterozygous positive factor V Leiden mutation | 1344 | 1344 | Factual
follow-up MRV | 1344 | 1344 | Factual
complete recanalization of the thrombosed sinuses | 1344 | 1344 | Factual
no new thrombi | 1344 | 1344 | Factual
complete remission | 1680 | 1680 | Factual
regular follow-up | 1680 | 1680 | Factual
no other thrombotic events | 1680 | 1680 | Factual
no leukemia relapses | 1680 | 1680 | Factual