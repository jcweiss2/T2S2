39 years old | 0
female | 0
chronic kidney disease | -79200
maintenance hemodialysis | -79200
severe pulmonary artery hypertension | -79200
chronic pulmonary thromboembolism | -79200
progressive breathlessness | -168
abdominal distension | -168
Grade III dyspnea | 0
orthopnea | 0
no fever | 0
no cough | 0
blood pressure 92/46 mmHg | 0
pulse rate 96/min | 0
respiratory rate 36/min | 0
recurrent hypotension | -96
non-tolerance to hemodialysis | 0
peritoneal dialysis planned | 0
severe hypotension | 0
altered sensorium | 0
shifted to ICU | 0
drowsy | 0
sluggishly responding to verbal commands | 0
distended neck veins | 0
respiratory distress | 0
active accessory muscles of respiration | 0
loud P2 | 0
pan systolic murmur | 0
soft abdomen | 0
mildly distended abdomen | 0
free fluid | 0
palpable liver | 0
blood pressure 70/40 mmHg | 0
pulse rate 102/min | 0
respiratory rate 30/min | 0
SpO2 99% on high flow O2 | 0
hemoglobin 12.3 g/dl | 0
total leucocyte count 8600/μL | 0
serum sodium 138 mEq/L | 0
serum potassium 6 mEq/L | 0
blood urea nitrogen 63 mg/dl | 0
creatinine 6.0 mg/dl | 0
hypoxia | 0
hypercarbia | 0
mixed acidosis | 0
pH 7.189 | 0
PaCO2 60.3 mmHg | 0
pO2 52.7 mmHg | 0
HCO3 22.5 mmol/L | 0
BE 6.54 mmol/L | 0
serum lactate 1.92 mmol/L | 0
high D-dimer | 0
high fibrin degradation product | 0
dilated right ventricle | 0
dilated right atrial | 0
dilated inferior vena cava | 0
moderate tricuspid regurgitation | 0
severe pulmonary arterial hypertension | 0
PASP 93 mmHg | 0
paradoxical septal motion | 0
decreased right ventricular function | 0
reduced left ventricular compliance | 0
sepsis ruled out | 0
acute myocardial ischemia ruled out | 0
high dose inotropes | 0
vasopressors | 0
infusion nor-adrenaline 1 mcg/kg/min | 0
infusion dopamine 20 mcg/kg/min | 0
empiric broad spectrum antibiotics | 0
low molecular weight heparin | 0
sustained low efficiency dialysis | 0
increased vasopressor requirement | 24
infusion vasopressin 0.04 units/min | 24
poor sensorium | 24
hemodynamic instability | 24
acidosis | 24
elective intubation | 24
ventilation | 24
pre-intubation pH 7.18 | 24
pre-intubation PaCO2 60 mmHg | 24
pre-intubation PO2 66.6 mmHg | 24
pre-intubation HCO3 21.9 mmol/L | 24
pre-intubation BE 7.1 mmol/L | 24
post-intubation pH 7.29 | 24
post-intubation PaCO2 36.7 mmHg | 24
post-intubation PO2 80.4 mmHg | 24
post-intubation HCO3 17.3 mmol/L | 24
post-intubation BE 8.3 mmol/L | 24
echocardiography similar findings | 48
refractory pulmonary hypertension | 72
inhaled nitric oxide started | 72
nitric oxide blender | 72
iNO at 5 ppm | 72
iNO increased to 10 ppm | 72
improving hemodynamic parameters | 72
vasopressors tapered down | 84
peritoneal dialysis restarted | 120
cumulative negative balance 2 L | 120
pH 7.45 | 120
PaCO2 28.4 mmHg | 120
PO2 136.2 mmHg | 120
HCO3 20 mmol/L | 120
BE 5.3 mmol/L | 120
lactates 1.61 mmol/L | 120
PASP 73 mmHg | 120
PASP 63 mmHg | 144
vasopressors weaned off | 168
nitric oxide withdrawn | 168
extubated | 192
non-invasive ventilation | 192
inspiratory positive airway pressure 12 mmHg | 192
expiratory positive airway pressure 4 mmHg | 192
shifted out of ICU | 240
methemoglobin levels < 1% | 240
acute right heart syndrome | 0
chronic pulmonary artery hypertension decompensation | 0
multifactorial causes | 0
rescue treatment with inhaled nitric oxide | 72
acute management of hypoperfused state | 240
clinical improvement | 240
decrease in vasopressor requirement | 84
decrease in PASP | 120
successful weaning | 168
