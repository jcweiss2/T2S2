89 years old | 0
male | 0
admitted to the hospital | 0
vomiting | -96
epigastric distension | -96
no bowel movements | -96
no flatus | -96
gallstones | -8760
intermittent right upper quadrant pain | -8760
hypertension | 0
diabetes | 0
pulmonary tuberculosis | -43800
schistosomiasis | -43800
moderate drinking | 0
no smoking | 0
no allergies | 0
unremarkable family history | 0
temperature 36.2 °C | 0
heart rate 77 beats per min | 0
respiratory rate 20 breaths per min | 0
blood pressure 137/74 mmHg | 0
abdominal tenderness | 0
hyperactive bowel sounds | 0
normal lung examination | 0
normal heart examination | 0
normal routine blood examination | 0
normal liver function | 0
normal renal function | 0
normal coagulation function | 0
normal troponin | 0
normal procalcitonin | 0
high-sensitivity C-reactive protein increased | 0
abdominal contrast CT | 0
pneumatosis in the gallbladder | 0
cholecystoduodenal fistula | 0
gallstone in the upper jejunum | 0
intestinal obstruction | 0
pneumobilia | 0
Rigler’s triad | 0
magnetic resonance cholangiopancreatography | 0
short T2 signal | 0
intestinal dilatation | 0
propulsive enteroscopy | 24
deep ulcer in the duodenal bulb | 24
yellow purulent secretion | 24
mucosal edema | 24
stone incarceration | 24
food residue | 24
laser lithotripsy | 24
sodium bicarbonate injection | 24
second propulsive enteroscopy | 48
stone smaller | 48
laser lithotripsy | 48
sodium bicarbonate injection | 48
laparoscopic duodenoplasty | 192
cholecystectomy | 192
enterolithotomy | 192
repair | 192
severe inflammation | 192
edema around the gallbladder | 192
cholecystoduodenal fistula formation | 192
jejunal gallstone ileus | 192
gallbladder removal | 192
cauliflower drainage tube | 192
purse-string suturing | 192
jejunum cut | 192
gallstone removal | 192
intestine wall sutured | 192
drainage tubes | 192
tachycardia | 216
atrial fibrillation | 216
mild anemia | 216
hypoproteinemia | 216
elevated urea | 216
elevated creatinine | 216
elevated NT-proBNP | 216
deslanoside | 216
amiodarone hydrochloride | 216
sinus rhythm | 216
hypourocrinia | 240
anuria | 240
hyperpyrexia | 240
disturbance of consciousness | 240
elevated white blood cells | 240
coagulation abnormalities | 240
elevated troponin | 240
elevated NT-proBNP | 240
elevated creatinine | 240
elevated procalcitonin | 240
high-sensitivity C-reactive protein increased | 240
Enterococcus faecium | 240
meropenem | 240
tigecycline | 240
linezolid | 240
teicoplanin | 240
continuous renal replacement therapy | 240
intravenous plasma transfusion | 240
coronary dilating drugs | 240
abdominal tenderness | 264
rebound tenderness | 264
exudate around drainage tube | 264
hypotension | 264
noradrenaline | 264
pituitrin | 264
decrease in platelet count | 264
teicoplanin | 264
urine volume recovery | 288
stable vital signs | 288
decrease in white blood cell count | 432
moderate anemia | 432
elevated creatinine | 432
elevated troponin | 432
elevated NT-proBNP | 432
elevated procalcitonin | 432
cefoperzone sodium | 432
tazobactam sodium | 432
lethargy | 456
mouth breathing | 456
coma | 480
unresponsive pupils | 480
abdominal CT | 480
postoperative changes | 480
exudative effusion | 480
chest CT | 480
infection in the right lung | 480
head CT | 480
cerebral infarction | 480
anti-infective therapy | 480
supportive treatments | 480
enteral nutrition | 480
electrolytes maintenance | 480
oxygen therapy | 480
death | 504