42 years old | 0
    female | 0
    health care provider | 0
    presented to emergency department | 0
    high-grade fever | -48
    productive cough | -48
    shortness of breath | -48
    bony pains | -48
    history of contact with patient with similar complaints | -96
    left nephrectomy in 2012 for staghorn calculus | -336
    cesarean section 3 times | -336
    abortion once | -336
    obese | 0
    newly diagnosed with diabetes mellitus type 2 | 0
    not on diabetic medication | 0
    Glasgow Coma Scale 15/15 | 0
    hemodynamically stable | 0
    leukopenia | 0
    white cell count 3.7 | 0
    lymphopenia 0.39% | 0
    chest x-ray bilateral infiltrates | 0
    admitted to ward | 0
    septic screen for MERS-CoV | 0
    influenza AB test | 0
    H1N1 test | 0
    dengue serology | 0
    malaria test | 0
    started on broad spectrum antibiotics | 0
    started on oseltamivir | 0
    symptoms progressed | 0
    admitted to ICU | 0
    chest x-ray extensive bilateral consolidations | 0
    refractory hypoxemia | 0
    electively intubated | 0
    mechanically ventilated | 0
    100% Fraction of inspired oxygen | 0
    ARDS protocol | 0
    low tidal volume | 0
    prone position | 0
    tracheal aspirates sent for MERS-CoV PCR | 0
    MERS-CoV PCR positive | 0
    started on Peginterferon Alpha-2a | 0
    started on ribavirin | 0
    started on intravenous methylprednisolone 60 mg every 6 hours | 0
    extracorporeal membrane oxygenation contemplated | 0
    respiratory function improved | 120
    FiO2 40% | 288
    Partial Pressure of Oxygen 103.5 mm Hg | 288
    weaning trial planned | 288
    sedation cessation | 288
    methylprednisolone tapered to 40 mg IV every 6 hours | 288
    Peginterferon Alpha-2a discontinued | 288
    ribavirin discontinued | 288
    hemodynamically stable | 288
    respiratory function improved | 288
    chest consolidation improved | 288
    wake up | 288
    move all limbs | 288
    polyuria | 312
    urine osmolarity 95 | 312
    serum osmolarity 341 | 312
    urine sodium <20 | 312
    serum sodium 161 meq/L | 312
    chloride 119 meq/L | 312
    blood sugar 25 mmol/L | 312
    Desmopressin 2 ug subcutaneously | 312
    planned brain CT | 312
    unresponsive | 312
    GCS dropped to 3/15 | 312
    pupils 3 mm wide with sluggish reaction | 312
    CT brain right frontal hematoma | 312
    subarachnoid hemorrhage | 312
    intraventricular extension | 312
    midline shift | 312
    subfalcine herniation | 312
    normal platelet count 347 X 10^9 | 312
    normal coagulation profile | 312
    no anticoagulation treatment | 312
    blood cultures negative | 312
    intracranial bleed acute | 312
    intracranial bleed large | 312
    no surgical intervention | 312
    medical supportive measures | 312
    lost brain stem reflexes | 312
    pupils fixed and dilated | 312
    follow-up brain CT complete loss of gray and white matter differentiation | 312
    large frontal hematoma | 312
    complete effacement of extra axial CSF spaces | 312
    contrast-enhanced CT no vessel enhancement beyond internal carotid arteries | 312
    CT angiogram no visualization of Middle cerebral artery | 312
    no visualization of Posterior cerebral artery | 312
    no flow within posterior circulation | 312
    complete brain anoxia | 312
    lack of intracranial flow | 312
    brain death criteria | 312
    supportive measures continued | 312
    cardiac arrest | 2664
    declared dead | 2664
    <|eot_id|>
