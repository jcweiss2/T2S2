68 years old | 0
male | 0
admitted to the hospital | 0
history of coronary artery disease | 0
history of hypertension | 0
history of type II diabetes mellitus | 0
history of paroxysmal supraventricular tachycardia | 0
returned to the United States from the Philippines | 0
visited family in Manila | -2160
visited family in Lucena | -2160
developed myocardial infarction | -2160
hospitalized for myocardial infarction | -2160
received angioplasty | -2160
placement of two stents in coronary arteries | -2160
discharged from hospital in the Philippines | -1440
hospitalized for fevers and left upper quadrant abdominal pain | -720
discharged from hospital in the Philippines | -720
presented to the emergency room with progressive worsening of left upper quadrant abdominal pain | 0
temperature 97.5°F | 0
blood pressure 127/69 mmHg | 0
pulse 117 beats per minute | 0
respiration rate 27 breaths per minute | 0
oxygen saturation 99% on room air | 0
tenderness in the left upper quadrant on palpation | 0
CT scan of the abdomen and pelvis with intravenous contrast | 0
multiple ill-defined hypodense lesions in the spleen | 0
started empirically on oral ciprofloxacin and metronidazole | 0
changed to intravenous vancomycin, ceftazidime, and metronidazole | 0
blood cultures drawn prior to administration of antibiotics returned negative for growth | 0
urine culture returned positive for Group B streptococcus | 0
transthoracic echocardiogram performed | 0
no valvular vegetation or new regurgitant valvular pathology | 0
CT-guided aspiration of the splenic lesion | 48
culture of the aspirate grew Burkholderia pseudomallei | 48
antibiotic regimen changed to intravenous ceftazidime alone | 48
discharged on this regimen | 0
induction therapy with ceftazidime for 8 weeks | 0
eradication therapy with oral doxycycline and trimethoprim-sulfamethoxazole for 20 weeks | 0
complete resolution of fever, leukocytosis, and abdominal pain | 1680
repeat CT scan of the abdomen showed resolution of the splenic lesions | 1680
aspirate culture plate sent to the California Department of Public Health for confirmation of diagnosis | 0
diagnosis confirmed | 0
plate destroyed before antibiotic sensitivity testing could be performed | 0