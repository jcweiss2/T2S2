35 years old | 0
female | 0
resection of giant cell tumor | 0
right hand radius bone | 0
arthroplasty | 0
preoperative routine investigations | -24
coagulation profile | -24
standard monitors | 0
heart rate monitoring | 0
ECG monitoring | 0
noninvasive blood pressure monitoring | 0
pulse oximetry | 0
peripheral intravenous access |C0
supraclavicular brachial plexus block | 0
paresthesia technique | 0
anatomical landmarks | 0
third attempt | 0
paresthesia elicited | 0
0.5% bupivacaine | 0
2% lignocaine with adrenaline | 0
chest pain | 0
ipsilateral infraclavicular region | 0
chest expansion | 0
air entry | 0
X-ray chest | 0
no pneumothorax | 0
no fluid collection | 0
sedation with midazolam | 0
adequate sensory blockade | 0
adequate motor blockade | 0
surgery duration | 1.5
shifted to recovery room | 1.5
chest discomfort | 1.5
stable vitals | 1.5
heart rate 94/min | 1.5
respiratory rate 16/min | 1.5
blood pressure 119/68 mmHg | 1.5
SpO2 99% | 1.5
repeat chest X-ray | 1.5
oxygen supplementation | 1.5
sedation | 1.5
analgesia | 1.5
shifted to ward | 1.5
symptom free for 12–14 h | 14
chest pain | 14
palpitations | 14
reduced chest expansion | 14
absent air entry | 14
X-ray chest | 14
massive fluid collection | 14
partial lung collapse | 14
shifted to operation theater | 14
heart rate 119/min | 14
respiratory rate 30/min | 14
blood pressure 94/56 mmHg | 14
SpO2 96% | 14
oxygenation | 14
fluid resuscitation | 14
large-bore IV access | 14
intercostal tube drainage | 14
blood drainage 1300 ml | 14
blood cross-matching | 14
emergency investigations | 14
arterial gas analysis | 14
metabolic acidosis | 14
respiratory alkalosis | 14
hemothorax evacuation | 14
administered fresh whole blood | 14
shifted to ICU | 14
propped up position | 14
oxygen | 14
analgesics | 14
antibiotics | 14
ICU stay 5 days | 118
X-ray chest | 118
complete lung expansion | 118
retained hemothorax | 118
CT guided thoracoscopic evacuation | 118
discharged | 240
satisfactory condition | 240
