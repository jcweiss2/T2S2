66 years old | 0
    male | 0
    admitted to the hospital | 0
    10-day history of fever | -240
    fever | -240
    cough | -240
    sputum production | -240
    progressive jaundice | -240
    chronic alcoholic | -240
    drinking two or more bottles of liquor daily | -240
    diabetes mellitus | -240
    liver cirrhosis | -240
    cerebral infarction | -35040
    no neurological sequelae | -35040
    visited a hospital nearby | -240
    plain chest X-ray | -240
    abdominal computerized tomography (CT) scan | -240
    bilateral lower lung field haziness | -240
    27-mm liver mass | -240
    suspicion of aspiration pneumonia | -240
    suspicion of hepatocellular carcinoma | -240
    transferred to a secondary hospital | -240
    three days of intravenous antibiotics (ceftriaxone and azithromycin) | -72
    fever persisted | -72
    difficulty swallowing food | -72
    reflexive cough while drinking water | -72
    intact gag reflexes | 0
    decreased pharyngeal elevation | 0
    swollen bilateral anterior neck area | -336
    persisted for the last two weeks | -336
    lower left quadrant of the anterior neck swollen | -336
    mild tenderness | -336
    follow-up plain radiograph of the chest | 0
    normal chest radiograph | 0
    leukocytosis | 0
    WBC count: 18,690/µl | 0
    neutrophilia | 0
    89% of WBC | 0
    CRP increased to 14.8 mg/dl | 0
    VFSS performed | 0
    soft tissue posterior to the upper esophagus severely swollen | 0
    retropharyngeal mass | 0
    mechanical obstruction | 0
    laryngeal elevation restricted | 0
    epiglottic rotation restricted | 0
    aspiration occurred in all types of food | 0
    high risk of suffocation on puree-like diet | 0
    moderate-to-severe grade residues in the valleculae | 0
    moderate-to-severe grade residues in the pyriform sinuses | 0
    recommended tube feeding | 0
    nasogastric tube insertion unsuccessful | 0
    obstruction by the retropharyngeal mass | 0
    urgent contrast-enhanced CT scan of the neck | 0
    loculated fluid collection in the retropharyngeal space | 0
    loculated fluid collection in the anterior cervical space | 0
    loculated fluid collection in the pericarotid space | 0
    loculated fluid collection in the prevertebral space | 0
    fluid collection in the upper mediastinum | 0
    airway severely narrowed in the subglottic region | 0
    reactive intraparotid lymph nodes | 0
    reactive superficial cervical lymph nodes | 0
    left side of the neck | 0
    retropharyngeal abscess | 0
    mediastinitis | 0
    emergency tracheostomy | 24
    incision to drain the abscess | 24
    afebrile postoperative period | 24
    intravenous administration of ampicillin-sulbactam | 24
    culture of purulent discharge | 24
    methicillin-resistant Staphylococcus aureus | 24
    Klebsiella pneumoniae | 24
    administered ceftriaxone-vancomycin | 24
    CRP decreased to 10.2 mg/dl | 120
    transferred to the general ward | 240
    examination on the 18th postoperative day | 432
    general condition improved | 432
    follow-up VFSS performed | 432
    supraglottic penetration with curd-type yogurt | 432
    supraglottic penetration with large amount of free fluid | 432
    pharyngeal residue markedly reduced | 432
    recommended initiation of oral feeding training | 432
    nasogastric tube feeding maintained | 432
    tracheostomy tube removed | 504
    third VFSS performed | 648
    very little silent aspiration | 648
    teaspoon of fluid | 648
    recommended initiation of full oral feeding | 648
    puree-like consistency | 648
    follow-up chest CT | 648
    improvement in mediastinal extension | 648
    WBC count normalized to 7,510/µl | 648
    CRP normalized to 0.19 mg/dl | 648
    discharged | 1104
    swallowing function continued to improve | 1104
    stable full oral intake | 1104