62 years old | 0
male | 0
admitted to the hospital | 0
severe epigastric pain | -72
shortness of breath | -72
septic | 0
tachypnoeic | 0
tachycardic | 0
hypotensive | 0
temperature spiked to 38 °C | 0
blood sugar of 20 mmol/L | 0
intravenous insulin | 0
bilateral lung base crepitations | 0
distended abdomen | 0
crepitus in right lumbar region | 0
crepitus extending to scrotum | 0
rapid clinical deterioration | 0
cardiopulmonary resuscitation | 0
intubated | 0
inotropic support | 0
white cell count of 70 | 0
thrombocytopaenia of 14 | 0
C-reactive protein of 248 | 0
deranged renal profile | 0
serum creatinine of 578 | 0
urea of 47.6 | 0
coagulopathy | 0
mild transaminitis | 0
severe metabolic acidosis | 0
absence of the right kidney on ultrasonography | 0
gas production in the renal parenchyma | 0
air locules in anterior/posterior liver space | 0
air locules in retroperitoneum | 0
air locules in lateral abdominal muscle |C:\Users\b\AppData\Local\Temp\sumeplugins\plugins\outputFormatters\outputFormatterPy\f_3\62_yo_male_admitted_with_septic_shock_and_epn.txt
