53 years old | 0
male | 0
Caucasian | 0
admitted to hospital | 0
dyspnoea | -336
chest pain | -336
tachypnoea | 0
tachycardia | 0
elevated inflammatory markers | 0
CRP 105.8 mg/L | 0
multiple hospital attendances | -672
recurrent viral pericarditis | -672
non-steroidal anti-inflammatories | -672
colchicine | -672
prednisolone | -672
asthma | 0
allergic rhinitis | 0
hypertension | 0
hypercholesterolaemia | 0
obesity | 0
treated obstructive sleep apnoea | 0
afebrile | 0
normoxic | 0
normotensive | 0
tachycardic | 0
tachypnoeic | 0
soft dual heart sounds | 0
decreased breath sounds | 0
no pulsus paradoxus | 0
jugular venous pressure not elevated | 0
multiple previous fillings | 0
no over gingival inflammation | 0
no dental abscesses | 0
no decay | 0
sinus tachycardia | 0
no diffuse changes | 0
no electrical alternans | 0
normal white cell count | 0
elevated C-reactive protein | 0
chest X-ray unremarkable | 0
NTproBNP unremarkable | 0
autoimmune screens unremarkable | 0
mild left ventricular dysfunction | 0
large pericardial effusion | 0
organized echogenic material | 0
diastolic collapse | 0
significant tricuspid and mitral inflow variation | 0
dilated and fixed IVC | 0
pericardiocentesis | 0
150 mL blood-stained fluid drained | 0
symptom relief | 0
haemodynamic improvement | 0
pericardial fluid biochemistry | 0
lactate dehydrogenase 3584 U/L | 0
fluid/serum LD ratio 12 | 0
cholesterol concentration 1.7 mmol/L | 0
cultures sent | 0
pigtail catheter placed | 0
catheter removed | 48
minimal output | 48
improved inflammatory markers | 48
purulent debris observed | 48
repeat TTE | 48
small residual effusion | 48
RV free wall akinetic | 48
adherent | 48
ventricular interdependence | 48
minimally collapsing dilated IVC | 48
pericardial fluid cultured gram-positive bacillus | 48
i.v. vancomycin commenced | 48
targeted i.v. benzylpenicillin | 96
fungal and acid-fast bacilli cultures negative | 96
no malignant cells | 96
extensive workup negative | 96
repeat TTE | 96
increasing pericardial effusion | 96
worsening tricuspid and mitral inflow variation | 96
cardiac magnetic resonance imaging | 96
pericardial effusion | 96
markedly thickened pericardium | 96
constrictive effusive pericarditis | 96
no pulmonary infection | 96
surgical source control | 96
multidisciplinary meeting | 96
inpatient surgery | 120
significant exertional dyspnoea | 120
escalating inflammatory markers | 120
median sternotomy | 144
significant collection | 144
thickened pericardium | 144
purulent fluid drained | 144
pericardium resected | 144
right pleura opened | 144
drains inserted | 144
drains removed | 168
histopathology | 168
organizing fibrinous pericarditis | 168
reactive stromal and endothelial cells | 168
no malignant cells | 168
no bacterial growth | 168
surgical tissue acid-fast bacilli culture negative | 168
surgical tissue acid-fast bacilli microscopy negative | 168
blood, urine, and sputum cultures negative | 168
post-operative TTE | 168
small pericardial space | 168
no effusion | 168
preserved LV function | 168
discharged | 240
i.v. benzylpenicillin | 240
oral amoxicillin | 240
no further episodes | 720
low mood | 720
primary care physician | 720