75 years old | 0
man | 0
admitted to the cardiac care unit | 0
congestive heart failure | 0
non-ST elevated myocardial infarction | 0
CHF | 0
hypertension | 0
diabetes | 0
bronchial asthma | 0
hyperuricemia | 0
denied any past surgical interventions | 0
intubated | 0
underwent percutaneous coronary angioplasty | 0
refractory respiratory failure | 0
pulmonary edema | 0
pneumonia | 0
intubated three times in 18 days | 0
steroids | 0
intravenous methylprednisolone 40 mg | 0
switched to oral prednisone 30 mg | 72
tapering to 5 mg over 12 days | 72
ceftriaxone | 96
extubated on hospital day 18 | 432
routine chest radiography | 432
pneumomediastinum | 432
subcutaneous emphysema | 432
subdiaphragmatic free air | 432
afebrile | 432
vital signs normal | 432
mild tachycardia | 432
heart rate 105 bpm | 432
abdominal bloating | 432
denied abdominal pain | 432
crepitation all over his body | 432
abdomen distended | 432
abdomen soft | 432
white cell count 1.21x10^9/L | 432
blood urea nitrogen 89.6 mg/dL | 432
creatinine 4.35 mg/dL | 432
non-contrast CT | 432
subcutaneous emphysema over the chest and abdominal wall | 432
pneumomediastinum without pneumothorax | 432
massive pneumoperitoneum | 432
pneumoretroperitoneum | 432
diffuse mesenteric emphysema | 432
no ascites | 432
acute care surgery service consulted | 432
exploratory laparotomy | 432
gush of air evacuated | 432
no free fluid in the peritoneum | 432
diffuse emphysema in the small and large intestinal mesenteries and retroperitoneum | 432
mild emphysema and edema from the descending colon to the sigmoid colon | 432
no diverticula observed on the surface of the intestine | 432
examination of the intestine from stomach through rectum | 432
no perforation | 432
no discoloration | 432
descending colon not mobilized from the retroperitoneum | 432
abdomen closed | 432
transferred to the surgical intensive care unit | 432
extubated on postoperative day 1 | 456
transferred to the ward on postoperative day 2 | 480
postoperative day 9 | 576
fever spiked | 576
left lower quadrant pain | 576
septic shock | 576
blood specimens sent for culture | 576
sputum specimens sent for culture | 576
urine specimens sent for culture | 576
CT of the chest and abdomen with intravenous and oral contrast | 576
fat stranding | 576
extraluminal air | 576
small amount of free fluid around the descending colon | 576
returned to the operating room for re-exploration | 576
small abscess cavity identified in the mesentery of the descending colon | 576
Hartmann's procedure performed | 576
resected specimen | 576
tiny diverticulum penetrating the mesentery | 576
abscess formed | 576
pathological analysis compatible with perforated diverticulitis | 576
postoperative course complicated with prolonged mechanical ventilation | 576
tracheostomy | 576
discharged to a rehabilitation hospital | 1656
