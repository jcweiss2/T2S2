16 years old | 0
male | 0
Jamaican | 0
admitted to the hospital | 0
fatigue | -2160
epistaxis | -2160
dyspnea | -2160
white cell count of 1900 per cubic millimeter | -2160
absolute neutrophil count 90 per cubic millimeter | -2160
hemoglobin 5.3 g per deciliter | -2160
platelets 36 000 per cubic millimeter | -2160
hospitalized | -2160
bone marrow biopsy | -96
aplastic anemia | -96
discharged | -96
received packed red blood cells | -96
pooled platelet transfusions | -96
intravenous antibiotics | -96
admitted to the US National Institute of Health Clinical Center | 0
fever | -168
dysphagia | -168
odynophagia | -168
cough | -168
scant hemoptysis | -168
body temperature 38.2oC | 0
blood pressure 126/91 mm Hg | 0
heart rate 88 beats per minute | 0
respiratory rate 18 breaths per minute | 0
oxygen saturation 98% | 0
thin | 0
lethargic | 0
spitting blood-tinged saliva | 0
denies dyspnea | 0
phonating normally | 0
tender diffusely around the neck | 0
white cell count of 1430 per cubic millimeter | 0
absolute neutrophil count 0 per cubic millimeter | 0
hemoglobin 10.7 g per deciliter | 0
platelets 33 000 per cubic millimeter | 0
radiographic imaging showed a classic “thumbprint” sign | 0
direct laryngoscopy showed an erythematous, enlarged, and posteriorly ptotic epiglottis | 0
intravenous piperacillin/tazobactam | 0
vancomycin | 0
micafungin | 0
intravenous dexamethasone | 0
nebulized racemic epinephrine | 0
clinically improved | 24
blood cultures showed no growth | 24
endoscopically directed cultures from directly observed exudate on the right tonsillar area isolated Enterobacter cloacae | 24
prescribed meropenem | 24
follow-up laryngoscopy showed significant improvement | 408
discharged | 408