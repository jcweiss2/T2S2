66 years old | 0
    man | 0
    presented | 0
    intermittent high-grade fever | -2160
    generalized dullBcering abdominal pain | -2160
    passing turbid urine | -240
    decrease in urine output | -240
    swelling of both feet | -240
    treated with intravenous medications | -168
    type II diabetes mellitus | -26208
    regular medication for diabetes | -26208
    conscious | 0
    afebrile | 0
    tachycardic | 0
    heart rate of 136/min | 0
    blood pressure 110/70 mmHg | 0
    renal angle tenderness bilaterally | 0
    high total leukocyte counts | 0
    left shift | 0
    elevated urea | 0
    elevated creatinine | 0
    pyuria | 0
    leukocyte esterase positivity | 0
    possibility of pyelonephritis | 0
    possibility of renal abscess | 0
    acute kidney injury | 0
    activated partial thromboplastin time prolonged | 0
    sepsisBinduced coagulopathy | 0
    enlarged kidneys | 0
    bilateral renal abscesses | 0
    emergency ultrasoundBguided drainage of renal abscesses | 0
    transfusion of blood products | 0
    pus smear for bacterial culture | 0
    pus smear for fungal culture | 0
    pus smear for mycobacterial culture | 0
    GenExpert polymerase chain reaction test for Mycobacterium tuberculosis | 0
    X-ray chest normal | 0
    electrocardiogram normal | 0
    initiated on intravenous meropenem | 0
    adjusted for renal impairment | 0
    septate fungal hyphae | 0
    advised intravenous voriconazole | 0
    opted for intravenous amphotericin B | 0
    amphotericin B 1 mg/kg/day | 0
    Aspergillus fumigatus growth | 0
    worsening renal function | 0
    acute pulmonary edema | 0
    hyperkalemia | 0
    metabolic acidosis | 0
    initiated on hemodialysis | 0
    initiated on noninvasive ventilation | 0
    sudden cardiac arrest | 216
    aspiration | 216
    succumbed to illness | 216
    <|eot_id|>
    