20 years old | 0
    female | 0
    admitted to the hospital | 0
    dyspnea | -24
    cough | -72
    yellow sputum | -72
    intermittent fever | -72
    night sweats | -72
    exposure to upper respiratory infection | -168
    exposure to family member with recent travel to Morocco | -168
    visited buffalo farm | -168
    ate unpasteurized cheese | -168
    diffuse bilateral opacities on chest X-ray | 0
    severe hypoxemia | 0
    antibiotics initiated | 0
    admitted to ICU | 0
    community acquired pneumonia diagnosis | 0
    denied GI symptoms | 0
    denied rash | 0
    denied arthralgia | 0
    denied thromboembolic disease | 0
    denied chest pain | 0
    denied leg pain | 0
    denied swelling | 0
    oral contraceptive use | 0
    non-invasive positive pressure ventilation failure | 72
    intubation | 72
    echocardiogram showing normal cardiac function | 72
    respiratory cultures negative | 72
    enterovirus/rhinovirus detected | 72
    high PEEP | 72
    low tidal volume ventilation | 72
    hypoxemia (PaO2/FiO2 = 75) | 72
    hypercapnia | 72
    dense bilateral opacities with central air bronchograms | 72
    ECMO initiated | 72
    vancomycin | 0
    piperacillin-tazobactam | 0
    levofloxacin | 0
    high-dose intravenous vitamin C initiated | 72
    chest X-ray improvement | 96
    hemodynamic instability | 72
    vasopressor requirements | 72
    careful fluid balance management | 72
    bronchoscopy negative for pathogens | 120
    negative Histoplasma | 120
    negative Blastomyces | 120
    negative Aspergillus | 120
    negative Legionella antigen | 120
    furosemide use | 72
    daily negative fluid balance | 72
    continued resolution of lung opacities | 96
    improved lung gas exchange | 96
    further reduction in lung opacities | 168
    ECMO decannulation | 168
    extubation | 168
    vitamin C dosing reduced by half | 168
    vitamin C dosing reduced again by half | 192
    post-extubation requiring 4 L/min nasal oxygen | 168
    discharged home on room air | 288
    follow-up chest X-ray at 2 weeks post-discharge | 720
    completely recovered at 1 month follow-up | 720
    