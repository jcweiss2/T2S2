19 years old | 0  
    male | 0  
    admitted to the hospital | 0  
    persistent fever | -168  
    body ache | -168  
    throat pain | -168  
    decreased oral intake | -168  
    low blood pressure (systolic 90 mmHg) | 0  
    low blood pressure (diastolic 40 mmHg) | 0  
    normal saline infusion (1500 ml) | 0  
    shifted to medical intensive care unit | 0  
    broad-spectrum antibiotic started | 0  
    inotropic support (noradrenaline) started | 0  
    dengue test negative | 0  
    typhoid test negative | 0  
    malaria test negative | 0  
    leptospira test negative | 0  
    deranged kidney function tests | 0  
    deranged liver function tests | 0  
    pancytopenia | 0  
    coagulation disturbance | 0  
    hepatosplenomegaly | 0  
    HLH suspected | 0  
    laboratory investigations for HLH | 0  
    bone marrow biopsy performed | 0  
    intubated | 0  
    IV methylprednisolone pulse started | 0  
    TPE started | 0  
    elevated lactate dehydrogenase (2860 IU/L) | 0  
    low fibrinogen (50 mg/dl) | 0  
    elevated ferritin (3210 ng/ml) | 0  
    elevated fasting triglyceride (619 mg/dl) | 0  
    hemophagocytosis in bone marrow | 0  
    TPE sessions (3 consecutive days) | 72  
    IV dexamethasone maintenance started | 72  
    blood transfusion (2 units packed red cells) | 0  
    FFP transfusion (18 units) | 0  
    single donor platelet concentrates (4 units) | 0  
    cryoprecipitate transfusion (24 units) | 0  
    extubated | 72  
    discharged | 384  
    Hb 11.6 g/dl | 72  
    absolute neutrophil count 3.62 ×109/L | 72  
    platelet count 98 ×109/L | 72  
    PT/INR 13.5 | 72  
    fibrinogen 152 mg/dl | 72  
    fasting triglyceride 245 mg/dl | 72  
    serum ferritin 250 ng/ml | 72  
    improved organ function | 72  
    hematological parameters normalized | 384  
    biochemical parameters normalized | 384  
    coagulation parameters normalized | 384  

