47 years old | 0
female | 0
obese | 0
BMI of 42 | 0
admitted to the hospital | 0
incisional hernia | 0
hypertension | -672
transabdominal gynecologic surgery | -672
peripheral vascular disease | -672
angioplasties of the iliac arteries | -672
carbon dioxide pneumoperitoneum | 0
intraabdominal pressure 12mm Hg | 0
laparoscopic correction | 0
adhesiolysis | 0
15-minute break | 120
decompression of the abdomen | 120
pneumoperitoneum 215 minutes | 0
blood pressure stable | 0
hernia defect 20 cm × 16 cm | 0
expanded polytetrafluoroethylene meshes | 0
tackers | 0
transabdominal sutures | 0
paralytic ileus | 72
distended bowel | 72
C-reactive protein raised | 72
relaparoscopy | 72
intraabdominal pressure 12 mm Hg | 72
bowel distension | 72
no signs of contamination | 72
no signs of perforation | 72
no signs of ischemia | 72
systemic inflammatory response syndrome | 96
respiratory insufficiency | 96
transfer to intensive care unit | 96
bloody diarrhea | 216
colonoscopy | 216
severe ischemic colitis | 216
mesenteric angiography | 216
occluded superior mesenteric artery | 216
compensatory distended inferior mesenteric artery | 216
pinpoint stenosis | 216
balloon angioplasty | 216
anticoagulants | 216
improved | 216
deteriorated | 264
colonoscopy | 264
multiple perforations | 264
ischemic transverse colon | 264
laparotomy | 264
fecal peritonitis | 264
multiple perforations | 264
ischemic ascending and transverse colon | 264
resection of ischemic colon | 264
contaminated meshes removed | 264
deteriorated | 288
died | 288
histological examination | 288
extensive ischemia | 288
transmural ulcerations | 288
perforations | 288