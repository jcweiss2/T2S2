30 years old | 0
female | 0
admitted to the hospital | 0
abnormal liver function | -8760
persistent jaundice | -720
abdominal distension | -720
intermittent mild fever | -720
serologic antibodies negative | 0
antibodies of autoimmune diseases negative | 0
alpha fetoprotein negative | 0
no alcohol abuse | 0
no hepatotoxic prescriptions | 0
no gastrointestinal hemorrhage | 0
no surgery | 0
abdominal contrast-enhanced CT | -168
liver cirrhosis | -168
moderate ascites | -168
no space occupying lesions | -168
temperature 38.1°C | 0
heart rate 98 bpm | 0
normal breathing | 0
normal blood pressure | 0
fully conscious | 0
thyroid non-tender | 0
no thyromegaly | 0
bulging abdomen | 0
positive ascites sign | 0
pitting edema | 0
ecchymosis | 0
total leukocyte count 3.19 × 10^9/L | 0
neutrophil percentage 63.3% | 0
red blood cell count 3.46 × 10^12/L | 0
hemoglobin 10.7 g/L | 0
platelets 80 × 10^9/L | 0
bone marrow biopsy normal | 0
no infection | 0
liver function worsened | 0
increasing bilirubin | 0
coagulopathy | 0
low serum ceruloplasmin | 0
high urinary copper | 0
normal blood copper | 0
Kayser Fleischer ring | 0
positive gene detection of ATP-7B | 0
Wilson disease | 0
thyroid-stimulating hormone <0.005 mU/L | 0
free thyroxine 50.67 pmol/L | 0
thyrotrophin receptor antibody 4.52 IU/L | 0
Doppler ultrasound of thyroid abnormal | 0
anti-thyroid drugs contraindicated | 0
radioactive iodine therapy considered | 0
iodine level in 24-h thyroid uptake low | 0
anti-copper treatment not effective | 0
liver transplantation considered | 0
adjuvant medications used | 0
persistent mild fever | 0
liver function deteriorated | 0
hepatic encephalopathy | 384
coma | 432
plasma exchange | 432
mechanical ventilation | 432
supportive treatments | 432
persistently comatose | 432
increasing serum bilirubin | 432
bleeding in gastrointestinal | 432
bleeding in respiratory | 432
bleeding in urinary tract | 432
treatment stopped | 432
died | 432