51 years old | 0
    male | 0
    hypertension | 0
    admitted | 0
    pyogenic spondylodiscitis | 0
    severe COVID-19 illness | -336
    mechanical ventilation | -336
    ventilator-associated pneumonia | -336
    carbapenem-resistant Acinetobacter baumannii | -336
    ampicillin-sulbactam | -336
    polymyxin B | -336
    central line-related bloodstream infection | -336
    carbapenem-resistant Pseudomonas aeruginosa | -336
    meropenem | -336
    sacral pressure injury | -336
    critical illness polyneuropathy/myopathy | -336
    hospitalized for 57 days | -336
    hospital discharge | -672
    insidious pain in the lumbar region | -672
    insidious pain in the right hip | -672
    progressive worsening pain | -672
    impaired ambulation | -672
    no fever | -672
    no sphincter symptoms | -672
    severe pain on palpation of the lumbar spine | 0
    severe pain on mobilization of the lumbar spine | 0
    moderate pain in the right hip | 0
    normal muscle strength | 0
    normal reflexes | 0
    normal sensitivity | 0
    hemoglobin level of 12.1 g/dL | 0
    total leukocyte count of 8700 cells/mm³ | 0
    erythrocyte sedimentation rate of 120 mm/hr | 0
    C-reactive protein level of 1.5 mg/dL | 0
    computed tomography of the right hip | 0
    periarticular calcifications | 0
    heterotopic ossifications | 0
    magnetic resonance imaging of the lumbar spine | 0
    bone edema in T12 and L1 vertebral bodies | 0
    irregularity of the vertebral endplate | 0
    involvement of the psoas muscles | 0
    T12-L1 spondylodiscitis | 0
    psoitis | 0
    negative blood cultures | 0
    CT-guided bone biopsy | 48
    microbiological culture | 48
    Pseudomonas aeruginosa | 48
    susceptible to polymyxin B | 48
    susceptible to ceftazidime$avibactam | 48
    resistant to meropenem | 48
    resistant to imipenem | 48
    resistant to cefepime | 48
    resistant to ceftazidime | 48
    resistant to ciprofloxacin | 48
    resistant to piperacillin$tazobactam | 48
    resistant to tigecycline | 48
    resistant to amikacin | 48
    initiation of polymyxin B | 672
    initiation of meropenem | 672
    widespread cutaneous rash | 912
    switched to ceftazidime$avibactam | 912
    dermatological lesions disappeared | 912
    improvement in inflammatory markers | 912
    improvement in pain | 912
    tolerance to rehabilitation exercises | 912
    no adverse events | 912
    seven weeks of antimicrobial treatment | 1344
    conservative treatment for heterotopic calcification | 1344
    nonsteroidal anti-inflammatory drugs | 1344
    physical therapy | 1344
    improvement of hip pain | 1344
    complete return to work | 1824
    asymptomatic | 1824
    negative inflammatory markers | 1824
    healing of the spondylodiscitis | 1824
    resolution of bone edema | 1824
    absence of intervertebral or paravertebral fluid | 1824
    spondylodiscitis cure | 1824
    <|eot_id|>
    