54 years old | 0
male | 0
admitted to the hospital | 0
fevers | -120
vomiting | -120
non-productive cough | -120
shortness of breath | -120
lethargy | -120
collapsing | -120
left shoulder swelling | -120
left elbow redness | -336
chronic shoulder pain | -8760
bilateral shoulder dislocations | -8760
right humeral arthrodesis | -8760
alcohol misuse | -8760
paracetamol | -720
ibuprofen | -720
Kussmaul breathing | 0
heart rate of 115 | 0
blood pressure of 178/105 | 0
respiratory rate of 32 | 0
oxygen saturations of 98% | 0
elevated body mass index (BMI) of 30 | 0
increased work of breathing | 0
left renal angle tenderness | 0
warm erythematous and fluctuant swelling to his left elbow | 0
purulent draining sinus in his left axilla | 0
bedside glucose of 18.7 mmol/L | 0
ketones of 0.5 mmol/L | 0
acute kidney injury (AKI) | 0
urea of 10.1 mmol/L | 0
creatinine of 186 mmol/L | 0
thrombocytosis | 0
leukocytosis | 0
CRP of 424 mg/L | 0
deranged liver function tests (LFTs) | 0
elevated INR of 1.9 | 0
mixed metabolic acidosis | 0
hyperchloremic metabolic acidosis | 0
partial respiratory compensation | 0
anion gap of 20 mmol/L | 0
hypoalbuminaemia | 0
low serum potassium | 0
pyroglutamic acidosis suspected | 0
IV n-acetylcysteine (NAC) | 0
IV sodium bicarbonate | 0
liberal potassium supplementation | 0
peripherally inserted central catheter (PICC) | 0
computed tomography (CT) of his left upper limb and abdomen/pelvis | 12
collections in the left elbow, biceps and shoulder | 12
left-sided pyelonephritis | 12
incision, drainage and washout of his multiple collections | 24
MSSA bacteraemia | 24
disseminated infection | 24
cutaneous tissues of the left shoulder, left kidney, left inguinal lymph nodes and lungs | 24
transthoracic and transoesophageal echocardiogram | 24
non-invasive ventilation (NIV) for type 1 respiratory failure | 48
metastatic staphylococcal pneumonia | 48
IV cefazolin | 48
flucloxacillin sensitive | 48
elevated PGA level of 9 mmol/mmol of creatinine | 168
metformin | 168
gliclazide | 168
T2DM | 168
discharged | 672
representation to hospital | 720
delayed wound healing | 720
conservative management | 720