22 years old| 0
male| 0
presented to a primary care hospital with pain | -48
presented to a primary care hospital with tightness in the left upper abdomen | -48
presented to a primary care hospital with shortness of breath | -48
pain | -48
tightness in the left upper abdomen | -48
shortness of breath | -48
repeated episodes of mild to moderate breathlessness | -variable (past history)
consulted local physicians | -variable (past history)
prescribed symptomatic treatment | -variable (past history)
air fluid level in the left hemithorax | -48
diagnosed as hydropneumothorax | -48
left-sided intercostal drain (ICD) inserted | -48
serosanguinous fluid drained | -48
intercostal drains not relieved symptoms | -variable
second ICD inserted | -variable (after first ICD)
fluid stained with blood drained | -variable (after first ICD)
temporary relief of respiratory symptoms for a day | -24
low-grade fever | -24
pleuritic chest pain | -24
referred to our hospital | 0
unable to pass stool | -48
unable to pass flatus | -48
episodes of non-bilious vomiting | -48
febrile | 0
hemodynamically stable | 0
left ICDs in left hemithorax draining turbid foul-smelling contents | 0
decreased air entry on left lung | 0
abdominal viscera in left hemithorax | 0
fluid in left hemithorax | 0
abdominal tenderness | 0
guarding | 0
rigidity | 0
moderate respiratory embarrassment | 0
use of intercostal muscles of respiration | 0
subphrenic recession | 0
absent bowel sounds | 0
pulse rate 122 per min | 0
blood pressure 90 mm Hg systolic | 0
blood pressure improved to 110/80 mm Hg | 0
respiratory rate 34–36 per min | 0
pulse oximetry saturation 92–94% | 0
mild hypoxemia (paO2 72 mm Hg) | 0
mild metabolic acidosis (pH 7.31) | 0
serum bicarbonate 18 mmoles/liter | 0
air-fluid level in left hemithorax | 0
two ICDs in situ | 0
signs of peritonitis | 0
signs of sepsis | 0
emergency exploratory laparotomy | 0
general anesthesia induced | 0
crash induction performed | 0
ketamine 2 mg/kg | 0
fentanyl | 0
succinyl choline | 0
intubated with cuffed oral endotracheal tube | 0
oxygen | 0
nitrous oxide | 0
isoflurane | 0
vecuronium bromide | 0
intravenous fluids | 0
lactated ringers | 0
dextrose infused | 0
diaphragmatic defect (20×10 sq cm) | 0
stomach herniated into left chest | 0
splenic flexure of the colon herniated into left chest | 0
spleen herniated into left chest | 0
no peritoneal sac over stomach | 0
ICDs traumatized spleen | 0
ICDs traumatized stomach | 0
draining blood | 0
draining gastric contents | 0
tubes disconnected | 0
tubes removed | 0
splenectomy | 0
hernial contents reduced | 0
stomach perforation closed | 0
ICD placed in pleural cavity | 0
diaphragmatic defect repaired | 0
transfusion of two units packed red blood cells | 0
shifted to ICU | 0
respiratory support | 0
hemodynamic support | 0
neuromuscular blockade not reversed | 0
mild pleural effusion in left hemithorax | 0
lung re-expansion over three to five days | variable (postoperative days 3-5)
no lung hypoplasia | 0
extubated on fifth postoperative day | 120
hemodynamically stable postoperative course | variable (postoperative days)
chest expansion techniques | variable (postoperative)
physiotherapy | variable (postoperative)
transferred to general ward on seventh postoperative day | 168
recovered without further complications | variable
22 years old|0
male|0
presented to a primary care hospital with pain|-48
presented to a primary care hospital with tightness in the left upper abdomen|-48
presented to a primary care hospital with shortness of breath|-48
pain|-48
tightness in the left upper abdomen|-48
shortness of breath|-48
repeated episodes of mild to moderate breathlessness|-
consulted local physicians|-
prescribed symptomatic treatment|-
air fluid level in the left hemithorax|-48
diagnosed as hydropneumothorax|-48
left-sided intercostal drain (ICD) inserted|-48
serosanguinous fluid drained|-48
intercostal drains not relieved symptoms|-24
second ICD inserted|-24
fluid stained with blood drained|-24
temporary relief of respiratory symptoms for a day|-24
low-grade fever|-24
pleuritic chest pain|-24
referred to our hospital|0
unable to pass stool|-48
unable to pass flatus|-48
episodes of non-bilious vomiting|-48
febrile|0
hemodynamically stable|0
left ICDs in left hemithorax draining turbid foul-smelling contents|0
decreased air entry on left lung|0
abdominal viscera in left hemithorax|0
fluid in left hemithorax|0
abdominal tenderness|0
guarding|0
rigidity|0
moderate respiratory embarrassment|0
use of intercostal muscles of respiration|0
subphrenic recession|0
absent bowel sounds|0
pulse rate 122 per min|0
blood pressure 90 mm Hg systolic|0
blood pressure improved to 110/80 mm Hg|0
respiratory rate 34–36 per min|0
pulse oximetry saturation 92–94%|0
mild hypoxemia (paO2 72 mm Hg)|0
mild metabolic acidosis (pH 7.31)|0
serum bicarbonate 18 mmoles/liter|0
air-fluid level in left hemithorax|0
two ICDs in situ|0
signs of peritonitis|0
signs of sepsis|0
emergency exploratory laparotomy|0
general anesthesia induced|0
crash induction performed|0
ketamine 2 mg/kg|0
fentanyl|0
succinyl choline|0
intubated with cuffed oral endotracheal tube|0
oxygen|0
nitrous oxide|0
isoflurane|0
vecuronium bromide|0
intravenous fluids|0
lactated ringers|0
dextrose infused|0
diaphragmatic defect (20×10 sq cm)|0
stomach herniated into left chest|0
splenic flexure of the colon herniated into left chest|0
spleen herniated into left chest|0
no peritoneal sac over stomach|0
ICDs traumatized spleen|0
ICDs traumatized stomach|0
draining blood|0
draining gastric contents|0
tubes disconnected|0
tubes removed|0
splenectomy|0
hernial contents reduced|0
stomach perforation closed|0
ICD placed in pleural cavity|0
diaphragmatic defect repaired|0
transfusion of two units packed red blood cells|0
shifted to ICU|0
respiratory support|0
hemodynamic support|0
neuromuscular blockade not reversed|0
mild pleural effusion in left hemithorax|0
lung re-expansion over three to five days|72
no lung hypoplasia|0
extubated on fifth postoperative day|120
hemodynamically stable postoperative course|120
chest expansion techniques|120
physiotherapy|120
transferred to general ward on seventh postoperative day|168
recovered without further complications|168
