25 years old | 0
female | 0
low back pain | -72
intravenous drug use | -672
hypotension | -24
hypoxemic respiratory failure | -24
intubation | -24
tricuspid vegetations | -24
severe tricuspid regurgitation | -24
bilateral patchy opacifications | -24
pulseless electrical activity | -24
veno-arterial extracorporeal membrane oxygenation (VA-ECMO) | -24
norepinephrine | -24
methicillin-sensitive Staphylococcus aureus (MSSA) | 0
mildly reduced biventricular systolic function | 0
multiple tricuspid valve vegetations | 0
valve perforation | 0
severe tricuspid regurgitation | 0
lung consolidative and cavitary opacities | 0
small pleural effusions | 0
sacroiliitis | 0
no intracranial process | 0
differential hypoxemia | 24
conversion to VAV-ECMO | 24
percutaneous aspiration of tricuspid valve vegetations | 48
transition to VV-ECMO | 168
hypoxemia on VV-ECMO | 168
recirculation | 168
shunting of deoxygenated blood | 168
membrane dysfunction | 168
esmolol infusion | 240
reduction of cardiac output | 240
membrane lung shunting | 240
bronchopleural fistula | 336
empyema necessitans | 336
video-assisted thorascopic surgery | 336
Eloesser flap | 336
decannulation from VV-ECMO | 720
preserved left ventricular function | 720
dilated right ventricle | 720
normal systolic function | 720
persistent severe tricuspid regurgitation | 720
small vegetation | 720
discharge | 1440
no dyspnea | 4320
no symptoms of heart failure | 4320