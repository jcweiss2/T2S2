64 years old | 0
gentleman | 0
referred to the hospital | 0
acute pancreatitis | 0
Imrie/Glassgow Score = 6 | 0
biliary pathology | 0
initial CT scan of the abdomen | 0
extensive edematous changes involving the entire pancreas | 0
significant volume of HPVG | 0
concern regarding one segment of small bowel | 0
CT mesenteric angiogram | 2
poorly enhancing segment of small bowel | 2
venous thrombosis | 2
significant reduction in the volume of HPVG | 2
clinical condition disimproved | 2
emergency laparotomy | 2
resection of a nonviable ischemic segment of small bowel (60 cm) | 2
omental saponification | 2
prolonged intensive care admission (45 days) | 0
multiorgan dysfunction | 0
acute kidney injury | 0
adult respiratory distress syndrome | 0
discharged to the ward | 1080
readmitted to the intensive care unit | 1080 + 72 = 1152
overwhelming sepsis | 1152
repeat imaging | 1152
large peripancreatic necrotic collections | 1152
interventional radiology drainages | 1152
escalation in antimicrobials | 1152
escalation in antifungal | 1152
escalation in inotropic support | 1152
clinical condition deteriorated | 1152
died | 62 * 24 = 1488
male | 0
admitted to the hospital | 0
Imrie/Glasgow Score = 6 | 0
readmitted to the intensive care unit | 1152
died | 1488
