open modified Scopinaro procedure | -22896
weight reganance | -120
incisional hernia | -120
bariatric revisional surgery and hernia repair | -48
gastric pouch leak | -24
sepsis | -24
multiple intra-abdominal collections | -24
conservative management with open abdomen | -24
negative wound pressure therapy | -24
parenteral nutrition | -24
intravenous antibiotics | -24
epithelized gastrocutaneous fistula | -12
controlled but persistent drainage | -12
upper endoscopy | -12
fistulous orifice at the proximal edge of the vertical staple line | -12
extraluminal extravasation | -12
recurrent left subphrenic abscess | -12
endoscopic treatment | -12
argon plasma coagulation | -6
internal and external drainages | -6
clipping | -6
fibrin sealants | -6
e-vac therapy | -6
stenting | -6
multidisciplinary team discussion | 0
decision to proceed with an innovative endoscopic technique | 0
placement of a CSDO across the fistula orifice | 0
informed consent | 0
Occlutech® muscular VSD occluder placement | 2
intravenous sedation | 2
topic anesthesia | 2
fistula cannulation | 2
contrast injection | 2
AmplatzTM extra stiff guidewire insertion | 2
delivery system introduction | 2
CSDO deployment | 2
contrast study | 4
restricted oral intake | 24
liquid diet | 240
regular diet | 288
pigtail displacement | 1008
systemic signs of sepsis | 1008
computed tomography | 1008
fluoroscopy | 1008
partial dislodgment of the 8-mm mVSD CSDO | 1008
second attempt with an oversized disc | 1056
Occlutech® Figulla Flex II UNI 24-mm placement | 1056
upper endoscopy | 4320
contrast-enhanced CT scan | 4320
device engrafted | 4320
significant reduction of the chronic abscess | 4320
no signs of fistula recurrence | 4320
pigtail removal | 4320
no drainage | 4320