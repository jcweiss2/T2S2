76 years old | 0
male | 0
Caucasian | 0
admitted to the hospital | 0
hypertension | 0
type two diabetes mellitus | 0
stage four chronic kidney disease | 0
obstructive sleep apnoea | 0
previous pacemaker insertion | 0
previous bilateral total knee joint replacement | 0
chest pain | -48
shortness of breath | -336
electrocardiogram showed an old left bundle branch block | -48
high-sensitivity troponin levels 55 ng/L | -48
high-sensitivity troponin levels 71 ng/L | -46
temperature 35.8°C | -48
transthoracic echocardiography showed normal biventricular size and function | -48
angiography | -48
99% stenosis in a dominant right coronary artery | -48
four drug-eluting stents in the RCA | -48
balloon rupture | -48
discharged home | -72
represented with progressive shortness of breath | -24
mild bilateral pedal oedema | -24
normal heart and lung sounds | -24
white cell count of 14.3 × 10^9/L | -24
C-reactive protein of 110 mg/L | -24
non-dynamic high-sensitivity troponin levels of 85 ng/L | -24
non-dynamic high-sensitivity troponin levels of 82 ng/L | -24
transthoracic echocardiography showed normal biventricular function | -24
normal valve function with no evidence of endocarditis | -24
no pericardial effusion | -24
blood cultures positive | -16
started on IV flucloxacillin | -16
mild trauma to his left knee | -20
left knee aspirate | -12
left knee arthroscopic washout | -10
transoesophageal echocardiogram showed no evidence of endocarditis | -10
no pacemaker wire infection | -10
no pericardial effusion | -10
worsening shortness of breath | -8
pleuritic chest pain | -8
worsening kidney injury | -8
oliguria | -8
attempted dialysis | -6
hypotension | -6
angina | -6
admitted to intensive care unit | -4
dialysis with inotropic support | -4
focused cardiac ultrasound showed moderate pericardial effusion | -4
pericardiocentesis | -2
purulent pericardial fluid | -2
severe cardiogenic and vasoplegic shock | -2
hypoxia | -2
intubated | -2
computed tomography coronary angiography showed RCA aneurysm | 0
TTE showed severe biventricular failure | 0
large pericardial effusion | 0
pericardial drain blocks | 2
extubated | 6
percutaneous balloon pericardial window | 10
discharged from ICU | 14
discharged from hospital | 20
repeat TTE showed moderate to severely reduced left ventricular function | 720
moderately reduced right ventricular function | 720
no significant pericardial effusion | 720