61 years old | 0
woman | 0
presented to our hospital with pain in her right knee | 0
received a diagnosis of PJI after revision TKA | 0
given intravenous antibiotic treatment at the previous hospital | 0
referred to our hospital for treatment of septic shock | -24
had undergone primary TKA (Sigma RP-F, Depuy, Warsaw, IN, USA) for rheumatoid arthritis 10 years previously | -87600
revision TKA (P. F. C Sigma TC3, Depuy, Warsaw, IN, USA) due to aseptic loosening 6 months previously | -4320
receiving oral prednisone (4 mg daily) | -4320
tacrolimus (1.5 mg daily) | -4320
etanercept (50 mg subcutaneous injections weekly) | -4320
pain in the right knee | 0
swelling in the right knee | 0
burning sensations in the right knee | 0
redness in the right lower leg | 0
local heat in the right lower leg | 0
white blood cell count of 8.1×109/L | 0
C-reactive protein level of 19.9 mg/L | 0
aspiration of the right knee joint | 0
gram-positive streptococci detected by staining | 0
Streptococcus dysgalactiae (group G Streptococcus) identified | 0
temperature of 38.2°C | 0
heart rate of 128 beats/min | 0
blood pressure of 56/32 mmHg | 0
hemoglobin of 9.5 g/dL | 0
serum glucose of 99 mg/dL | 0
serum creatinine of 2.93 mg/dL | 0
sodium of 139 mEq/L | 0
radiography of the right knee showed no osteolytic lesions | 0
radiography of the right knee showed no signs of periprosthetic loosening | 0
computed tomography scan not performed | 0
diagnosed septic shock due to PJI after revision TKA | 0
rapidly performed irrigation | 0
debridement | 0
polyethylene liner exchange | 0
antibiotic therapy | 0
lack of tissue resistance to blunt finger dissection observed during surgery | 0
admitted to the Intensive Care Unit for mechanical ventilation | 0
placed empirically on meropenem (1.0 g every 12 h) | 0
vancomycin (0.5 g every 12 h) | 0
clindamycin (600 mg every 8 h) | 0
administered continuous hemodiafiltration | 0
started on nor-adrenaline via a peripheral intravenous catheter | 0
blood culture tests performed several times | 0
blood culture results all negative | 0
clinical condition gradually stabilized | 0
noradrenaline application stopped on day 5 of admission | 120
swelling in the right knee observed on hospitalization day 8 | 192
burning sensation in the right knee observed on hospitalization day 8 | 192
approximately 35 mL of exudate aspirated | 192
joint aspiration revealed white blood cell count of 60 100/ μL | 192
positive alpha-defensin test | 192
judged eradication failure of the infection | 192
performed irrigation | 192
debridement | 192
implant removal | 192
antibiotic spacer placement | 192
postoperative period was uneventful | 192
six weeks after surgery, inflammatory markers had normalized | 1008
intravenous antibiotic therapy (ampicillin 2 g every 6 h and clindamycin 600 mg every 8 h for 2 weeks) | 1008
cefazolin 2 g every 8 h for 4 weeks | 1008
ten weeks after surgery, no clinical signs of infection | 1680
discharged from the hospital with 2 canes | 1680
started on bucillamine (100 mg daily) 1 month after surgery | 720
dose gradually increased to 300 mg daily | 720
taking busiramine at discharge | 1680
taking prednisolone (4 mg daily) at discharge | 1680
bDMARDs not resumed | 1680
RA well controlled | 1680
administrated oral cefalexin 500 mg 3 times a day for 2 months | 1680
approximately 1.5 years after surgery, underwent re-revision TKA | 13104
inflammatory markers not elevated throughout the follow-up period | 13104
no clinical signs of infection observed throughout the follow-up period | 13104
one year after the final surgery, walked with a cane | 26208
no symptoms of infection | 26208
no pain in the right knee | 26208
no swelling in the right knee | 26208
no burning sensation in the right knee | 26208
right knee motion ranged from 0° of extension to 90° of flexion | 26208
no extension lag | 26208
