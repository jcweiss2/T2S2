62 years old | 0  
    male | 0  
    COVID-19 | -48  
    dyspnea | -48  
    asthenia | -48  
    fever (38°C) | -48  
    oxygen saturation (SaO2) of 93% | -48  
    cough | -48  
    hypertension | 0  
    left hydronephrosis (II-III grade) | 0  
    kidney stones | 0  
    bilateral pneumonia | 0  
    diffuse ground-glass opacity (GGO) | 0  
    clinical condition worsened | 0  
    admitted to ICU | 0  
    nasal intermittent positive pressure ventilation (NIPPV) | 0  
    Venturi mask with oxygen at 14 l/m | 0  
    pO2 of 42.5 mmHg | 0  
    pCO2 of 32.9 mmHg | 0  
    continuous positive airway pressure (CPAP) | 0  
    endotracheal intubation | 24  
    mechanical ventilation | 24  
    lung-protective ventilation with low-medium tidal volume (VT) at 6 mL/kg | 24  
    prone positioning | 24  
    Klebsiella pneumoniae infection | 336  
    consolidation in left lower lobe | 336  
    SaO2 stable above 90% | 336  
    D-dimer increased to 974 ng/mL | 336  
    Staphylococcus capitis infection | 504  
    Stenotrophomonas maltophilia infection | 504  
    bronchoaspiration | 504  
    severe hypoxemia | 504  
    ventilator maladjustment | 504  
    severe respiratory acidosis | 504  
    hypotension | 504  
    mechanical ventilation via tracheostomy | 720  
    death | 888  
    sepsis | 888  
    suppurative pericarditis | 888  
    mural thrombi in large heart vessels | 888  
    superficial microhemorrhagic areas in kidneys | 888  
    parenchymal congestion in kidneys | 888  
    necrotic area in liver | 888  
    liver parenchymal congestion | 888  
    glomerular collapse | 888  
    acute tubulointerstitial nephritis | 888  
    occasional renal arterioles thrombosis | 888  
    hepatic centrilobular vein thrombosis | 888  
    periportal inflammation | 888  
    hepatic sinusoids dilatation | 888  
    hepatic sinusoids congestion | 888  
    mild cholestasis | 888  
    increased lung parenchymal density | 888  
    whitish fibrotic areas in lungs | 888  
    pulmonary infarction areas | 888  
    advanced DAD | 888  
    collagen/fibrotic replacement tissue | 888  
    large protein globules | 888  
    vascular microthrombosis | 888  
    fibrosis with lumen obliteration | 888  
    fibroblasts present | 888  
    macrophages present | 888  
    type II hyperplastic pneumocytes present | 888  
    ventilator-induced lung injury (VILI) | 504  
    ventilator-associated lung injury (VALI) | 504  
    nosocomial bacterial superinfections | 504  
    polymicrobial lung superinfection | 504  
    pulmonary fibrosis | 888  
    cytokine activation | 888  
    multi-organ dysfunction syndrome (MODS) | 888  
    thromboembolism | 888  
    hypercoagulability | 888  
    mixed infections | 504  
    septic shock risk | 504  
    biofilm-related infections | 504  
    methicillin resistance | 504  
    pulmonary gangrene | 888  
    endotymological investigation lacking | 0  
    rapid bacterial infection detection | 0  
    patient isolation measures | 0  
    antimicrobial therapy management | 0  
    epidemiological monitoring | 0  
    family information provision | 0  