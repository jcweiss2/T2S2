18 years old | 0
male | 0
admitted to the hospital | 0
posterior uveitis | -168
testicular pain | -720
benign hypo-echoic lesions | -720
massive bleeding from mouth | 0
cardiac arrest | 0
cardiopulmonary resuscitation | 0
intubated | 0
ventilated | 0
shifted to intensive care unit | 0
endotracheal tube and nasogastric tube continued to drain over 500 ml of bloody aspirate | 0
esophagogastrodudenoscopy | 24
coffee ground material in stomach | 24
no signs of active bleeding | 24
toxicology screening negative | 24
autoimmune profile negative | 24
viral & Brucella serology negative | 24
Glasgow coma scale of 7 | 24
CT scan chest with contrast negative for pulmonary embolism | 24
echocardiogram suspicious for probable mass versus vegetation over tricuspid valve | 48
IV antibiotics | 48
antifungal | 48
second echocardiography | 72
cardiac surgery review | 72
discontinued all antibiotics/antifungal | 336
CT brain revealed hypoxic brain injury with minimal cerebral edema | 72
myoclonic seizures | 72
treated with phenytoin | 72
maintained on sodium valproate | 72
urologist’s impression that the lesions are likely secondary to a traumatic cause | 168
recurrent oral and genital ulcers | -720
recurrent joint pains | -720
Pathergy test inconclusive | 168
ophthalmological examination significant for posterior uveitis | 168
rheumatologist’s opinion | 168
treated with steroids | 168
CT chest with contrast showed massive pulmonary arteriovenous malformations/aneurysm | 168
left small pulmonary infarct | 168
Methylprednisolone 1 gram intravenous pulse therapy | 168
initiation of azathioprine 50mg | 168
steroids tapered down over 6 months | 720
maintained on 10 mg prednisolone with azathiprine 75 mg daily | 720
osteoporosis prevention medications | 720
extubated | 720
tracheostomy closed | 720
irreversible brain hypoxic injury | 720
minimal responsiveness with eye contact and nodding | 720
no motor response in the limbs | 720
follow-up with cardiology, rheumatology, nephrology and neurology | 720
biochemistry remained normal | 720
repeat ultrasound revealed that the testicular lesions had completely resolved | 876
repeat echocardiography revealed that the tricuspid lesion had also completely resolved | 876
repeat CT scan chest showed all pulmonary arterial aneurysms resolved | 876
discharged with home health care | 876
remained in an unchanged condition | 876
bedridden with persistent hypoxic brain injury | 876
no new lesions or other active problems | 876