21 years old | 0
male | 0
obese | 0
admitted to the hospital | 0
cough | -72
fever | -72
shortness of breath | -72
pleuritic chest pain | -72
light-headedness | -72
near syncope | -72
dyspnoea | -72
COVID-19 | 0
sub-massive pulmonary embolism | 0
unfractionated heparin | 0
hypotensive | 12
massive pulmonary embolism | 12
catheter-directed thrombolysis | 12
improved clinically | 24
discharge | 48
acute respiratory failure | 96
hypotension | 96
intubated | 96
cardiac arrest | 96
vasopressor support | 96
veno-arterial extracorporeal membrane oxygenation | 96
recurrent massive pulmonary embolism | 96
repeat catheter-directed thrombolysis | 96
ventilation parameters improved | 144
vasopressors discontinued | 144
venous duplex ultrasound | 144
deep venous thrombus | 144
inferior vena cava filter | 144
low-molecular-weight heparin | 144
pulmonary artery angiogram | 240
improvement in emboli burden | 240
weaned from ECMO | 240
decannulated | 240
septic shock | 336
broad spectrum antibiotics | 336
right thigh haematoma | 336
compartment syndrome | 336
surgical debridement | 336
rivaroxaban | 336
discharged | 1248
home | 2016
activities of daily living | 2016
anticoagulated | 2016
rivaroxaban | 2016