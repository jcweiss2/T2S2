67 years old | 0  
    Asian | 0  
    male | 0  
    attended the emergency room | 0  
    nausea | -24  
    vomiting | -24  
    diarrhoea | -24  
    fever | -24  
    lower abdominal pain | -24  
    no haematemesis | 0  
    no melena | 0  
    no urinary complaints | 0  
    passed eight watery bowel motions | 0  
    denied previous febrile illness | 0  
    denied sweating | 0  
    denied weight loss | 0  
    denied sexually transmitted disease | 0  
    past medical history unremarkable | 0  
    surgical history unremarkable | 0  
    drug history unremarkable | 0  
    no allergies | 0  
    businessman | 0  
    non-smoker | 0  
    no alcohol use | 0  
    performed Umrah | 0  
    looked sick | 0  
    dry mucous membranes | 0  
    temperature 38.7°C | 0  
    pulse rate 112/min regular | 0  
    blood pressure 140/90 | 0  
    oxygen saturation 98% | 0  
    severe tenderness at the right iliac fossa | 0  
    no rebound | 0  
    normal bowel sounds | 0  
    unremarkable heart exam | 0  
    unremarkable chest exam | 0  
    WBC count 24,000×109/l | 0  
    neutrophils 90% | 0  
    haemoglobin 10 g/dl | 0  
    normal MCV | 0  
    normal platelets | 0  
    serum creatinine 190 μmol/l | 0  
    urea nitrogen 12.5 mmol/l | 0  
    normal electrolytes | 0  
    normal liver function tests | 0  
    normal coagulation profile | 0  
    normal lactic acid | 0  
    stool analysis WBCs >20/hpf | 0  
    RBCs 3–5/hpf | 0  
    no ova | 0  
    no parasites | 0  
    negative blood culture | 72  
    negative stool culture | 72  
    negative Clostridium difficile PCR | 0  
    C-reactive protein 70 mg/l | 0  
    clinical picture suggesting acute gastroenteritis | 0  
    tenderness at the right iliac fossa | 0  
    received saline | 0  
    received paracetamol | 0  
    received ciprofloxacin 500 mg IV | 0  
    CT scan abdomen and pelvis without contrast | 0  
    AAA above renal arteries | 0  
    hyper-dense retroperitoneal haematoma | 0  
    intramural thrombus | 0  
    AAA 74 mm sagittal diameter | 0  
    aortic leak to right psoas muscle | 0  
    aortic leak to right iliac fossa | 0  
    good bilateral arterial pulsations | 0  
    transferred to vascular surgery team | 0  
    empirical antibiotics continued | 0  
    fever resolved | 0  
    inflammatory markers improved | 0  
    normal RPR serology | 0  
    normal chest x-ray | 0  
    exploratory laparotomy | 0  
    leaking juxtarenal AAA 10x7 cm | 0  
    aneurysm from renal artery to iliac bifurcation | 0  
    surgical repair | 0  
    intramural thrombus removed | 0  
    Dacron graft applied | 0  
    postoperative ICU admission | 0  
    received ventilation | 0  
    received inotropes | 0  
    correction of anaemia | 0  
    off ventilator after 2 days | 48  
    off inotropes after 2 days | 48  
    renal functions normalized by day 5 | 120  
    transferred to normal ward | 120  
    started rehabilitation | 120  
    discharged after 3 weeks | 504  
    flew back home | 504  
    ruptured AAA | 0  
    pain as presenting symptom | 0  
    abdominal pain | 0  
    flank/back pain | 0  
    hip pain | 0  
    testicular pain | 0  
    haematoma at left iliopsoas muscle | 0  
    left iliac fossa pain | 0  
    diarrhoea | 0  
    age as risk factor | 0  
    sex as risk factor | 0  
    acute bacterial gastroenteritis | 0  
    haematoma tracking to right iliac fossa | 0  
    intramural thrombus | 0  
    infectious AAA differential | 0  
    no previous febrile illness | 0  
    1-day gastroenteritis | -24  
    negative septic screen | 0  
    negative RPR | 0  
    hypotension | 0  
    shock related to sepsis | 0  
    adverse management outcome | 0  
   