30 years old | 0
female | 0
homozygous sickle cell disease | 0
admitted to the ICU | 0
respiratory failure | 0
neurological deterioration | 0
vaso-occlusive crisis | -72
fever | -72
pain in lower extremities | -72
lethargic | 0
temperature 38 ° | 0
heart rate 140 bpm | 0
anemia | 0
hemoglobin 8.3 g/dl | 0
decreased haptoglobin | 0
hyperleukocytosis | 0
PNN 18.7 × 10^3/μL | 0
CRP 215mg/L | 0
liver tests altered | 0
AST 121 UI/L | 0
ALT 64 UI/L | 0
AP 450 UI/L | 0
LDH 3861 UI/L | 0
total bilirubin 3.9 mg/dL | 0
renal function normal | 0
arterial oxygen saturation 80% | 0
chest CT angiography | 0
bilateral pulmonary consolidations | 0
pulmonary embolism excluded | 0
unenhanced cerebral CT-scan | 0
CT-angiography unremarkable | 0
SARS-CoV-2 RT-PCR negative | 0
SARS-CoV-2 serology negative | 0
diagnosis of vaso-occlusive crisis | 0
acute thoracic syndrome | 0
transferred to ICU | 0
MRI of the brain | 72
cerebral fat embolism syndrome | 72
punctate foci of restricted diffusion | 72
T2 FLAIR prolongation | 72
punctate foci of low signal intensity | 72
antalgics | 0
antibiotics | 0
red cell exchange | 0
discharged from ICU | 96
neurological symptoms regressed | 336
follow-up cerebral MRI | 8760
signal abnormalities regressed | 8760
cerebral microbleeds persistent | 8760