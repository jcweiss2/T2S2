44 years old | 0
woman | 0
right-sided facial paralysis | 0
removal of acoustic neuroma | 0
lagophthalmos | 0
continued keratopathy | 0
implantation of gold weight in right upper eyelid | 0
postoperative day 11 | 264
right eyelid swelling | 264
erythema | 264
limitation of abduction | 264
orbital cellulitis | 264
intravenous cefuroxime | 264
complete limitation of gaze | 264
afferent pupillary defect | 264
necrosis of lower eyelid | 264
necrosis of upper eyelid margins | 264
necrosis of anterior ocular segment | 264
computed tomography scan | 264
swelling of superficial tissues | 264
removal of gold weight | 264
necrosis in upper eyelid tarsus | 264
necrosis in lower eyelid | 264
necrosis in limbus | 264
necrosis in conjunctiva | 264
opaque cornea | 264
dense cataract | 264
full thickness biopsy of eyelid | 264
necrotic conjunctiva | 264
necrotic skin | 264
diffuse acute inflammatory reaction | 264
gram-positive cocci | 264
Staphylococcus capitis | 264
intravenous vancomycin | 264
piperacillin/tazobactam | 264
stabilization | 264
light perception only visual acuity | 264
transcranial Doppler | 264
normal flow in ophthalmic arteries | 264
four days following gold weight removal | 336
fever 38°C | 336
chills | 336
tachycardia | 336
extreme restlessness | 336
systemic involvement | 336
thinning of sclera | 336
necrosis of sclera | 336
worsening of eyelid swelling | 336
worsening of eyelid necrosis | 336
axial computed tomography scan with contrast | 336
air bubbles under eyelid | 336
intraconal fat haziness | 336
infectious or inflammatory process | 336
evisceration | 336
debridement of necrotic tissue | 336
acute nonspecific necrotizing panophthalmitis | 336
gram-positive cocci | 336
Staphylococcus epidermidis | 336
Candida albicans | 336
Candida glabrata | 336
clindamycin | 336
voriconazole | 336
deterioration | 336
fever | 336
urinary retention | 336
desaturation | 336
acidosis | 336
admission to intensive care unit | 336
stabilization | 336
vancomycin | 336
meropenem | 336
fluconazole | 336
improvement | 336
stable ocular condition | 336
severe contracted socket | 336
a year later | 8760
admitted to plastic surgery ward | 8760
5-month-old nonhealing third-degree chemical burn of right anterior thigh | 8760
wound debridement under local anesthesia | 8760
lack of patient cooperation | 8760
complete debridement under general anesthesia | 8760
split thickness skin graft | 8760
negative pressure dressing | 8760
postoperative day 2 | 8760
torn negative pressure dressing | 8760
dressing change | 8760
partially taken skin graft | 8760
Sulfamylon wet-to-dry dressing | 8760
tenderness | 8760
itching | 8760
unrest | 8760
postoperative day 11 | 8760
full thickness third-degree burn | 8760
no signs of infection | 8760
debridement | 8760
partial thickness skin graft | 8760
postoperative day 1 | 8760
torn dressing | 8760
torn skin graft | 8760
third skin grafting | 8760
full length cast | 8760
protection | 8760
immobilization | 8760
self-induced damage | 8760
high suspicion of factitious disorder | 8760
psychiatric consult | 8760
diagnosis of factitious disorder could not be made | 8760
