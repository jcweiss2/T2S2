50 years old | 0
male | 0
Vietnamese | 0
admitted to the intensive care unit | 0
diffuse abdominal pain | -168
vomiting | -168
watery diarrhea | -168
fever | -168
productive cough | -168
bilateral pleuritic chest pain | -168
intermittent asthma | -6720
seizure disorder | -6720
heavy alcohol drinker | -6720
severe respiratory distress | 0
tachycardic | 0
afebrile | 0
hypoxic | 0
borderline hypotension | 0
blood pressure of 90/60 mm Hg | 0
diffuse rhonchi | 0
intubation | 0
mechanical ventilation | 0
leucopenia | 0
thrombocytopenia | 0
lactic acidosis | 0
severe transaminitis | 0
bilateral infiltrates | 0
intravenous fluids | 0
broad-spectrum antibiotics | 0
vancomycin | 0
piperacillin tazobactam | 0
oseltamivir | 0
azithromycin | 0
septic shock | 0
pneumonia | 0
acute respiratory distress syndrome | 24
piperacillin | 24
tazobactam | 24
azithromycin | 24
meropenem | 24
levofloxacin | 24
leptospirosis | 24
fiberoptic bronchoscopy | 24
bronchoalveolar lavage | 24
Klebsiella pneumoniae | 24
parainfluenza | 24
propofol | 0
fentanyl | 0
lorazepam | 0
dexmedetomidine | 96
severe agitation | 96
weaning attempts | 96
acute abdominal distension | 216
ileus | 216
abdominal pain | 216
non-bloody diarrhea | 216
dilated cecum | 216
abdominal x-ray | 216
abdominal CT | 216
toxic megacolon | 216
volvulus | 216
nasogastric tube | 216
rectal tube | 216
electrolytes replacement | 216
fluid replacement | 216
antibiotics | 216
infectious colitis | 216
Clostridium difficile infection | 216
C. difficile toxin A and B | 216
GDH antigen | 216
stool for ova | 216
parasite | 216
culture | 216
endoscopic decompressions | 264
surgery | 264
cecal perforation | 264
serosal tear | 264
side-to-side ileocolic anastomosis | 264
diversion loop ileostomy | 264
patchy transmural suppurative acute and chronic inflammation | 264
ulceration | 264
mucosal necrosis | 264
serositis | 264
fungal hyphae | 264
ischemic colitis | 264
perforation | 264
ACPO | 264
discharged | 1008
skilled nursing facility | 1008
jejunostomy tube feeding | 1008
tracheostomy | 1008