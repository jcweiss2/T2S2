43 years old | 0
woman | 0
gradually gained weight | -17520
leg edema | -17520
referred to a clinic | -17520
nephrotic syndrome | -17520
admitted to a hospital | -17520
minimal change nephrotic syndrome | -17520
steroid therapy | -17520
steroid pulse | -17520
daily oral prednisolone | -17520
high fever | -168
acute kidney injury | -168
admitted to our hospital | 0
drowsy | 0
blood pressure 121/93 mmHg | 0
pulse rate 80/min | 0
body temperature 36.8°C | 0
bilateral lower extremity edema | 0
no chest pain | 0
no abdominal tenderness | 0
CRP 48.93 mg/dL | 0
Alb 1.4 g/dL | 0
CK 2529 mg/dL | 0
CK-MB 196 mg/dL | 0
Cr 3.75 mg/dL | 0
troponin-T 14.19 ng/mL | 0
PCT 100.0 ng/mL | 0
marked proteinuria | 0
nephrotic syndrome | 0
ST-elevation on ECG | 0
pleural effusion | 0
no pulmonary congestion | 0
reduced wall motion of left ventricle | 0
ejection fraction 30% | 0
hypokinesis | 0
Takotsubo cardiomyopathy | 0
acute myocarditis | 0
no significant elevation in antibody titers | 0
Escherichia coli in blood culture | 0
sepsis due to Escherichia coli | 0
Meropenem | 0
Levofloxacin | 0
severe respiratory distress | 24
pulmonary congestion | 24
anuria | 24
non-invasive positive pressure ventilation | 24
continuous hemodiafiltration | 24
slight calcification in left ventricle | 120
myocarditis recovery | 240
respiratory status recovery | 240
AKI improvement | 336
stop dialytic therapy | 336
Warfarin | 336
remission of MCNS | 744
reduce prednisolone dose | 744
discharged | 912
widespread calcification | 1344
impaired cardiac function | 1344
EF 46% | 1344
wall motion impairment at apex | 1344
delayed enhancement on MRI | 1344
calcification persistent | 8760
cardiac function slight improvement | 8760
