47 years old | 0
male | 0
admitted to the hospital | 0
persistent severe headache | -1080
computed tomographic imaging of the head | 0
diffuse bleed in the subarachnoid space | 0
anterior communicating artery aneurysm | 0
chronic smoker | 0
nonalcoholic | 0
no known comorbid illness | 0
neurological deterioration | -12
flexor response to painful stimuli | -12
fresh bleed | -12
hydrocephalus | -12
external ventricular drain | -12
sensorium improved | -6
emergency surgery | -6
permanent clips | -6
ventriculoperitoneal shunt | -6
elective ventilation | 0
extubated | 24
neurologically well preserved | 24
Glasgow Coma Scale E3M6V5 | 24
fever | 48
hypotension | 48
deterioration in sensorium | 48
Glasgow Coma Scale E2M5V2 | 48
sepsis suspected | 48
resuscitated with fluids | 48
antibiotics | 48
elective ventilation | 48
noradrenaline infusion | 48
repeat DSA | 48
complete clipping of the aneurysm | 48
no evidence of vasospasm | 48
abdominal distension | 72
persisting fever | 72
ultrasound examination of the abdomen | 72
moderate ascites | 72
bilateral pleural effusion | 72
severe hypoalbuminemia | 72
intravenous albumin | 72
elevated lipase | 96
normal serum amylase | 96
normal calcium | 96
normal triglyceride levels | 96
CT abdomen | 96
edematous pancreas | 96
peripancreatic fat stranding | 96
conservative management | 96
antibiotics | 96
antipyretics | 96
total parental nutrition | 96
fluctuations in sensorium | 168
externalization of VP shunt | 168
improved neurologic status | 168
laboratory testing of ascitic fluid | 168
no signs of infection | 168
tracheostomized | 240
weaned from the ventilator | 240
Glasgow Coma Scale E4M6Vt | 240
enteral feedings initiated | 240
lipase level returned to baseline | 240
fever | 336
altered sensorium | 336
redness | 336
induration | 336
purulent discharge | 336
subcutaneous swelling | 336
Klebsiella | 336
septic shock | 336
died | 344