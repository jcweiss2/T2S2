72 years old|0
    male|0
    fever|-72
    chills|-72
    cough|-72
    chest pain|-72
    high leucocyte count (37100/mm3)|0
    right lung consolidation (chest radiograph)|0
    low blood pressure|0
    transferred to ICU|0
    pneumonia|0
    septic shock|0
    noradrenaline infusion started (0.1 mcg/kg/min via peripheral IV)|0
    IV cannula placed (dorsum of left hand)|0
    broad-spectrum antibiotics|0
    fluid resuscitation|0
    vasopressor support|0
    blood pressure stabilized|0
    vasopressor tapering after 2 hours|120
    CVC placement not attempted|120
    swelling (dorsum of left hand)|12
    purplish discoloration|12
    infusion stopped|12
    IV cannula removed|12
    new IV cannula placed (volar aspect of right forearm)|12
    NA infusion tapered off|16
    NA infusion stopped|16
    topical nitroglycerin 2% applied (every 4 hours)|12
    hand elevation|12
    phentolamine unavailable|0
    terbutaline unavailable|0
    heat application|12
    swelling and discoloration improvement|24
    skin texture near normal after 48 hours|48
    
    72 years old|0
    male|0
    fever|-72
    chills|-72
    cough|-72
    chest pain|-72
    high leucocyte count (37100/mm3)|0
    right lung consolidation (chest radiograph)|0
    low blood pressure|0
    transferred to ICU|0
    pneumonia|0
    septic shock|0
    noradrenaline infusion started (0.1 mcg/kg/min via peripheral IV)|0
    IV cannula placed (dorsum of left hand)|0
    broad-spectrum antibiotics|0
    fluid resuscitation|0
    vasopressor support|0
    blood pressure stabilized|0
    vasopressor tapering after 2 hours|120
    CVC placement not attempted|120
    swelling (dorsum of left hand)|12
    purplish discoloration|12
    infusion stopped|12
    IV cannula removed|12
    new IV cannula placed (volar aspect of right forearm)|12
    NA infusion tapered off|16
    NA infusion stopped|16
    topical nitroglycerin 2% applied (every 4 hours)|12
    hand elevation|12
    phentolamine unavailable|0
    terbutaline unavailable|0
    heat application|12
    swelling and discoloration improvement|24
    skin texture near normal after 48 hours|48