17 years old | 0
female | 0
admitted to the Emergency Department | 0
fever | -264
altered behavior | -264
abnormal body movement | -264
altered sensorium | -264
agitation | -264
suspiciousness | -264
aggression | -264
restlessness | -264
sleep disturbance | -264
violent behavior | -264
olanzapine prescribed | -264
phenytoin prescribed | -264
temperature 101°F | 0
blood pressure 130/70 mmHg | 0
tachycardia | 0
heart rate 117 beats/min | 0
tachypnea | 0
respiratory rate 20 breaths/min | 0
oxygen saturation 92% | 0
Glasgow Coma Scale 8/15 | 0
Antibody Prevalence in Epilepsy and Encephalopathy score 7 | 0
absence of nuchal rigidity | 0
bilateral mute plantar reflex | 0
cognitive function not assessable | 0
oxygen therapy started | 0
intravenous fluids started | 0
anticonvulsants started | 0
antibiotics started | 0
transferred to ICU | 0
CT scan of head normal | 0
MRI of brain normal | 0
CT scan of abdomen and pelvis normal | 0
lumbar puncture performed | 0
CSF analysis showed lymphocytic pleocytosis | 0
protein and glucose normal in CSF | 0
RT-PCR for HSV-1 and HSV-2 negative | 0
RT-PCR for Mycobacterium tuberculosis negative | 0
autoimmune encephalitis panel sent | 0
anti-NMDA receptor antibodies positive | 0
diagnosis of anti-NMDA receptor encephalitis confirmed | 0
methylprednisolone started | 0
intravenous immunoglobulins started | 0
condition did not improve | 120
ventilator-associated pneumonia developed | 120
rituximab not administered | 120
septic shock developed | 144
vasopressor therapy started | 144
intractable cardiac failure | 168
death | 168