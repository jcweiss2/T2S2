55 years old | 0
female | 0
smoker | 0
chronic obstructive pulmonary disease | 0
diabetes | 0
admitted to the emergency department | 0
worsening dyspnea | 0
respiratory distress | 0
tachypnea | 0
tachycardia | 0
wheezing | 0
decreased breath sounds in the left upper lung field | 0
pneumonia | 0
acute respiratory failure | 0
intravenous antibiotics | 0
fluid resuscitation | 0
noninvasive ventilatory support | 0
right upper quadrant pain | 0
high alkaline phosphate level | 0
abdominal ultrasonography | 0
enlarged liver | 0
multiple masses | 0
chest computed tomography | 0
abdomen computed tomography | 0
7-cm mass in the left upper lung lobe | 0
obstructive pneumonitis | 0
extensive bilateral mediastinal and left hilar, axillary, and supraclavicular lymphadenopathy | 0
multiple liver metastases | 0
histopathologic examination | 0
liver biopsy | 0
high-grade small cell neuroendocrine cancer | 0
magnetic resonance imaging of the brain | 0
normal brain findings | 0
extensive stage small cell lung cancer | 0
oliguria | 96
elevated creatinine | 96
elevated potassium | 96
sepsis-associated acute kidney injury | 96
increasing potassium | 96
increasing phosphorus | 96
increasing uric acid | 96
spontaneous tumor lysis syndrome | 96
fluid resuscitation | 96
phosphate binders | 96
allopurinol | 96
rasburicase | 96
renal function deterioration | 120
elevated creatinine | 120
oncology consultation | 120
nephrology consultation | 120
daily hemolysis | 144
palliative chemotherapy | 144
cisplatin | 144
etoposide | 144
dialysis dependent | 216