47 years old | 0
male | 0
presented with 1-week history of melaena | -168
passing 2 dark, tarry stools per day | -168
experienced 7 months of proximal muscle weakness | -5040
12 kg of weight loss | -5040
using a walking stick due to right hip pain | -1008
low energy fall from a bicycle 6 weeks prior | -1008
medical history of grade 1 pancreatic head neuroendocrine tumour | -52560
tumour staged as T3N1M0 | -52560
Ki-67 index of <2% | -52560
non-functional tumour | -52560
serum chromogranin A normal | -52560
serum chromogranin B normal | -52560
gut hormone levels normal | -52560
underwent pylorus-preserving pancreaticoduodenectomy | -52560
on pancreatin | -52560
insulin glargine at night | -52560
insulin aspart with meals | -52560
sinus tachycardia of 115 beats per minute | 0
blood pressure 128/63 mm Hg | 0
bilateral pitting oedema to mid-thigh | 0
soft abdomen | 0
non-tender abdomen | 0
no hepatosplenomegaly | 0
digital rectal examination confirmed melaena | 0
haemoglobin 85 g/L | 0
acute drop from haemoglobin 120 g/L | -240
mildly raised urea 8.3 mmol/L | 0
normal creatinine 77 μmol/L | 0
hypokalaemic 2.9 mmol/L | 0
normal liver function | 0
normal coagulation profile | 0
normal albumin 41 g/L | 0
negative transthoracic echocardiogram | 0
negative oesophago-gastro-duodenoscopies | 0
negative colonoscopy | 0
negative video capsule endoscopy | 0
CT scan showing portal hypertension | 0
variceal dilatation of mesenteric veins | 0
no parenchymal liver disease | 0
no ascites | 0
no pleural effusions | 0
sub-acute right pubic rami fractures | -1008
gallium-68 DOTATATE PET showing SMV recurrence | 0
intraluminal SMV tumour invasion | 0
porto-mesenteric hypertension | 0
bleeding mesenteric varices | 0
managed conservatively with blood transfusions | 0
potassium replacement | 0
commenced on lanreotide autogel 120 mg monthly | 0
discharged after 24 days | 576
admitted to intensive care with septic shock | 672
Escherichia coli bacteraemia | 672
cytomegalovirus viraemia | 672
discharged to rehabilitation after 5 weeks | 1344
bedbound due to deconditioning | 1344
worsening proximal myopathy | 1416
lower back pain | 1416
unexplained ecchymosis | 1416
re-admitted to hospital | 1416
hypertensive 162/107 mm Hg | 1416
unexplained oedema | 1416
hypokalaemia 2.9 mmol/L | 1416
hypernatraemia 148 mmol/L | 1416
metabolic alkalosis pH 7.53 | 1416
bicarbonate 38.6 mmol/L | 1416
osteoporotic vertebral compression fractures | 1416
24-h urinary free cortisol collection | 1416
low-dose dexamethasone test | 1416
confirmed Cushing's syndrome | 1416
elevated ACTH levels | 1416
ectopic ACTH source | 1416
negative pituitary MRI | 1416
repeat gallium-68 DOTATATE PET scan | 1416
ectopic ACTH release from pNET recurrence | 1416
commenced on metyrapone 1000 mg TID | 1416
ketoconazole 200 mg TID | 1416
hydrocortisone 10 mg BID | 1416
normalized serum cortisol | 1416
discharged home after 27 days | 1944
continued lanreotide therapy | 1944
reduction in tumour size | 1944
community physiotherapy | 1944
regained near pre-morbid performance status | 1944
plans for chemotherapy | 1944
surgical resection deemed high risk | 1944
