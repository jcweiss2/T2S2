51 years old | 0
male | 0
white | 0
admitted to the hospital | 0
history of severe alcoholism | -8760
high daily consumption of alcohol | -8760
consumed rum | -8760
consumed cognac | -8760
consumed wines | -8760
refused to treat addiction | -8760
decrease in short-term memory | -876
paresthesias of the lower limbs | -876
paresthesias of the upper limbs | -876
ingestion of large amounts of alcohol | -24
excessive drowsiness | -24
torpor | -12
coma | 0
Glasgow coma score 7 | 0
no signs of meningeal irritation | 0
no focal deficits | 0
no cranial nerve abnormalities | 0
IV thiamine administration | 0
high doses of parenteral B vitamins administration | 0
hypodensity in the corpus callosum on CT scan | 0
involvement of the cortical regions and subcortical white matter on MRI | 0
mild improvement in level of consciousness | 24
Glasgow coma score 10 | 24
mechanical ventilatory support | 24
multiple pulmonary infectious complications | 168
respiratory insufficiency | 168
dependent on mechanical ventilation | 168
tracheostomy | 168
septic | 720
fever | 720
worsening of respiratory status | 720
hemodynamic condition deteriorated | 720
vasoactive drugs administration | 720
broad-spectrum IV antibiotics administration | 720
cultures of blood and tracheal secretions revealed Rhodotorula mucilaginosa | 720
amphotericin B treatment | 720
no significant response to amphotericin B | 744
septic shock | 744
death | 744