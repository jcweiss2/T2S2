54 years old | 0
woman | 0
admitted to hospital | 0
allergic reaction to amoxicillin | -6
single dose of amoxicillin | -6
suspected upper respiratory tract infection | -6
transient episodes of turning pale | -12960
transient episodes of feeling lightheaded | -12960
'white outs' | -12960
diffuse non-blanching rash | -6
blood pressure 192/122 mm Hg | -6
no clinical signs of airways obstruction | -6
chest tightness | 0
no wheeze | 0
no stridor | 0
diffuse mottled vasculitic rash (livedo reticularis) | 0
pyrexial | 0
hypertensive | 0
persistently tachycardic | 0
normal chest X ray | 0
elevated white cell count | 0
elevated C reactive protein | 0
deranged liver function | 0
deranged coagulation profile | 0
acute kidney injury | 0
treated for anaphylactic reaction to amoxicillin | 0
treated for systemic infection | 0
started on broad spectrum antibiotics | 0
started on intravenous fluids | 0
started on supportive therapy in intensive care unit | 0
became restless | 72
became agitated | 72
altered level of consciousness | 72
clinical features suggestive of global encephalopathy | 72
unremarkable CT head | 72
unremarkable lumbar puncture | 72
unremarkable initial septic screen | 72
atrial fibrillation | 72
fast ventricular rate | 72
drop in blood pressure | 72
received noradrenaline | 72
blood pressure remained labile | 72
discontinued noradrenaline after 72 h | 72
10 cm heterogeneous right adrenal mass on CT | 72
diagnosis of pheochromocytoma crisis considered | 72
given intravenous phentolamine | 72
confirmed pheochromocytoma crisis | 72
blood pressure stabilized within 36 h of phentolamine | 72
switched to oral phenoxybenzamine after four days | 96
cardiac arrest | 240
45 minutes of CPR | 240
ejection fraction 40% | 240
multi-organ failure | 240
low Glasgow Coma Scale | 240
continued to deteriorate | 384
died | 384
