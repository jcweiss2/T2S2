23 years old | 0
man | 0
presented with retrosternal pleuritic chest pain | 0
low-grade fever | 0
apyretic | 0
normotensive | 0
pericardial rub present | 0
electrocardiogram showed sinus tachycardia | 0
widespread ST elevation | 0
PR segment depression | 0
echocardiography showed mild circumferential pericardial effusion | 0
normal high sensitivity troponin I | 0
mild leukocytosis | 0
very elevated C-reactive protein | 0
developed cardiac tamponade | 24
emergent pericardiocentesis performed | 24
evacuation of 350 ml serous fluid | 24
progressed to profound shock | 24
dependent on high noradrenaline doses | 24
1-g bolus methylprednisolone administered | 24
excellent clinical response verified | 24
weaning of noradrenaline | 48
progressive resolution of effusion | 48
childhood asthma | -10080
nonallergic rhinitis | -10080
idiopathic episcleritis | -10080
controlled with topical corticosteroids | -10080
admitted to intensive care unit | -720
septic shock | -720
tonsillitis | -720
pericardial friction rub | 0
differential diagnosis of acute pericarditis | 0
differential diagnosis of myocarditis | 0
differential diagnosis of pulmonary embolism | 0
differential diagnosis of pneumonia | 0
differential diagnosis of asthma exacerbation | 0
differential diagnosis of pneumothorax | 0
Streptococcus mitis isolated in pericardial fluid | 0
ceftriaxone initiated | 0
echocardiogram showed constrictive-effusive physiology | 0
autoimmunity workup pendent | 0
discharged on colchicine | 0
ibuprofen | 0
prednisolone | 0
working diagnosis of idiopathic acute pericarditis | 0
readmitted due to incessant pericarditis | 672
cardiac tamponade | 672
immediate pericardiocentesis | 672
pleuro-pericardial window performed | 672
pericardial biopsy obtained | 672
cardiac magnetic resonance showed diastolic paradoxical septal movement | 672
diffuse pericardial late gadolinium enhancement | 672
discharged with higher dose methylprednisolone | 672
symptoms recurred when corticosteroid dose lowered to <10 mg | 672
several readmissions | 672
hyperkalemia | 672
hyponatremia | 672
suspicion of adrenal insufficiency | 672
adrenocorticotropin levels very high | 672
cortisol under limit of detection | 672
diagnosis of Addison's disease | 672
hormonal replacement therapy with fludrocortisone | 672
prednisolone | 672
anti-intrinsic factor autoantibodies present | 672
primary hypogonadism found | 672
diagnosis of autoimmune polyglandular syndrome type 2 | 672
free T4/TSH normal | 672
γ interferon negative | 672
HIV serology negative | 672
cytomegalovirus IgM/IgG negative/positive | 672
Epstein Barr virus IgM/IgG negative/positive | 672
parvovirus IgM/IgG negative/positive | 672
herpes virus 1 IgM/IgG negative/positive | 672
herpes virus 2 IgM/IgG negative/negative | 672
Coxiella burnetti negative | 672
Borrelia burgdoferi IgM/IgG negative/negative | 672
Rickettsia conori IgG positive | 672
Treponema pallidum negative | 672
antinuclear antibodies positive | 672
anti-dsDNA antibodies negative | 672
anti-pANCA/c ANCA negative | 672
anti-SSA60, Sm, RNP, Scl70, JO negative | 672
rheumatoid factor negative | 672
septic shock complicating tonsillitis | -720
recurrent cardiac tamponade | 672
shock | 672
high-dose bolus corticosteroid reverted shock | 24
methylprednisolone maintenance contributed to clinical response | 24
impaired response to stressful event | 672
adrenal crisis | 672
high mortality | 672
primary AI | 672
Addison's disease | 672
mineralocorticoid insufficiency | 672
APS-2 | 672
recurrence of pericarditis | 672
corticosteroid dependence | 672
prednisolone successfully tapered to 5 mg q.d. | 672
new recurrence | 672
required higher doses | 672
Addisonian crisis | 672
life-threatening situation | 672
multiple clinical presentations | 672
diagnosis challenging | 672
pericardial tamponade as first presentation | 672
broader etiological study motivated | 672
