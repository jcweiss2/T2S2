85 years old | 0
Caucasian woman | 0
homemaker | 0
rheumatoid arthritis | 0
hyperlipidemia | 0
asthma | 0
cerebrovascular accident (CVA) | -1440
second dose of MODERNA COVID-19 vaccine | -48
generalized weakness | -48
muscle cramps | -48
loss of appetite | -48
first dose of MODERNA vaccine | -768
minor pain at the injection site | -768
weak | -48
could not stand up from the toilet seat | -48
stayed in bed except while using the bathroom with assistance | -48
lost appetite | -48
nausea | -48
urine color changing from dark brown to black | -48
weakness worsened | -24
abdominal cramps | -24
muscle cramps | -24
brought to the ER by ambulance | -24
clopidogrel | -1440
metoprolol | 0
nifedipine | 0
rosuvastatin | 0
telmisartan | 0
tofacitinib | 0
trazodone | -1440
stroke | -1440
professional physiotherapy once a week | 0
non-weight bearing exercises daily | 0
family history of autoimmune disease | 0
no tobacco or alcohol abuse | 0
never contracted COVID-19 | 0
no recent trauma or surgery | 0
no recent over-the-counter medications | 0
exhausted | 0
hypoactive bowel sounds | 0
generalized mild abdominal tenderness | 0
alert and oriented | 0
stable vital signs | 0
elevated serum creatinine | 0
elevated BUN | 0
decreased GFR | 0
low bicarbonate | 0
elevated AST | 0
elevated ALT | 0
elevated alkaline phosphatase | 0
elevated CPK | 0
elevated troponin | 0
urinalysis positive for blood | 0
negative RBCs | 0
elevated myoglobin | 0
non-contrast CT abdomen negative | 0
non-contrast CT head negative | 0
elevated aldolase | 0
hemolysis | 0
bicarbonate-rich IV fluids | 0
heart failure with preserved ejection fraction (HFpEF) exacerbation | 0
elevated pro-BNP | 0
ejection fraction 55-60% | 0
diastolic dysfunction | 0
progressively weaker | 0
could not lift/move hands or legs | 0
mentation decline | 0
confusion | 0
hallucinations | 0
3+ pitting edema | 0
chest CT consolidation right lower lobe | 0
chest CT consolidation left lower lobe | 0
ascites | 0
anasarca | 0
broad-spectrum IV antibiotics | 0
temporary dialysis catheter | 0
hemodialysis | 0
hypoxia from pleural effusion | 0
oliguria | 0
renal failure | 0
empiric glucocorticoids | 0
myositis | 0
CSF clear | 0
negative CSF cultures | 0
elevated CSF glucose | 0
elevated CSF total protein | 0
elevated myelin basic protein | 0
negative VDRL | 0
negative herpes I/II | 0
negative West Nile | 0
transferred to ICU | 0
bilevel positive airway pressure | 0
high-flow oxygen | 0
intubated | 0
ventilator support | 0
CPK remained elevated | 0
cardiac arrest | 0
hypoxic/anoxic brain injury | 0
palliative care consultation | 0
terminally extubated | 0
died | 24
