23 years old | 0
male | 0
T-cell precursor lymphoblastic leukemia | -35040
allogenic stem cell transplantation | -35040
disease relapse | -96
re-induction therapy | -96
local radiotherapy | -96
systemic chemotherapy | -96
nelarabine | -96
triple intrathecal chemotherapy | -96
complete disease remission | -96
consolidation chemotherapy | -72
second allogenic stem cell transplantation | -72
GvHD prophylaxis | -72
cyclosporine | -72
methotrexate | -72
mild oral mucositis | -72
headache | -72
moderate abdominal discomfort | -72
slightly elevated CRP | -72
hyperpotassemia | -72
cyclosporine dosage reduced | -72
initial improvement of symptoms | -72
recurrent hyperpotassemia | -24
SPS 15 mg orally | -24
progressive abdominal pain | 0
fever | 0
tachycardia | 0
normotensive | 0
peripheral oxygen saturation normal | 0
abdomen bloated | 0
no signs of peritonitis | 0
leukopenia | 0
neutropenia | 0
elevated CRP | 0
CT scan | 0
thickened gastric wall | 0
gastric pneumatosis | 0
air in hepatic portal vein system | 0
upper GI endoscopy | 0
generalized mucosal erythema | 0
intramucosal bleeding | 0
necrosis of gastric fundus and corpus | 0
exploratory laparotomy | 0
necrosis of gastric wall confirmed | 0
total gastrectomy | 0
esophago-jejunal anastomosis | 0
postoperative intensive care | 0
transferred to isolation ward | 0
total parenteral nutrition | 0
antibiotic therapy | 0
histopathology | 0
ischemic transmural necrosis | 0
purulent peritonitis | 0
kayexalate crystals | 0
no GvHD | 0
no Helicobacter pylori infection | 0
vital resection margins | 0
upper GI X-ray series | 168
normal passage | 168
no leakage | 168
fully recovered | 168
discharged | 720
