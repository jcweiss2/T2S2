46 years old | 0
male | 0
admitted to the hospital | 0
sepsis | 0
left hip periprosthetic infection | 0
increased pain in the left hip | -24
drainage of blood and purulence | -24
open wound | -24
no history of trauma | 0
no preceding fevers or chills | 0
psoriatic arthritis | -672
treated with steroids | -672
treated with methotrexate | -672
left metal-on-metal THA | -648
right metal-on-metal THA | -324
elevated white blood cell count | 0
decreased hemoglobin | 0
elevated C-reactive protein | 0
elevated erythrocyte sedimentation rate | 0
decreased albumin | 0
blood cultures drawn | 0
radiograph of the pelvis, left hip, and left femur | 0
hemodynamically stable | 0
no shortness of breath | 0
denies chest pain | 0
vancomycin | 0
Zosyn | 0
negative deep vein thrombosis ultrasound | 0
normal electrocardiogram | 0
physical examination | 0
temporal wasting | 0
severe bilateral lower extremity psoriasis | 0
no neurovascular deficits | 0
fungating mass | 0
left hip pain | -2592
radiographs of the pelvis and left hip | -2592
computed tomography of the abdomen and pelvis | -2592
mild particle wear | -2592
left hip fluid collection | -2592
aspiration | -2592
intravenous vancomycin | -2592
intravenous Zosyn | -2592
orthopaedic consultation | -2592
aspirated culture negative | -2592
antibiotics stopped | -2592
discharged | -2592
left hip pain | -1092
radiographs of the hip and pelvis | -1092
MRI | -1092
CT | -1092
loss of the left hemipelvis | -1092
bubbling osteolysis | -1092
massive pseudotumor | -1092
bone loss | -1092
acetabulum | -1092
hemipelvis | -1092
worked up for infection | -1092
worked up for metallosis | -1092
serum chromium | -1092
serum cobalt | -1092
elevated erythrocyte sedimentation rate | -1092
elevated C-reactive protein | -1092
aspiration | -1092
three-dimensional reconstruction CT scan | -1092
surgery | -1092
cup-cage construct | -1092
custom triflange | -1092
allograft hemipelvis reconstruction | -1092
aspiration results negative | -1092
no antibiotics | -1092
three-dimensional scans | -1092
DePuy Synthes | -1092
modeling of the pelvis | -1092
revision of failed left THA | -1092
metallosis | -1092
debridement of the pseudotumor | -1092
intraoperative biopsy | -1092
acute-on-chronic inflammation | -1092
cultures negative | -1092
intraoperative finding | -1092
bearing surface wear | -1092
intraoperative biopsy results | -1092
acute-on-chronic inflammation | -1092
cultures negative | -1092
discharged | -1092
follow-up | -1092
radiographs | -1092
continued erosion | -1092
left hemipelvis | -1092
proximal femur | -1092
left hip disarticulation | 48
surgical planning | 48
elevated inflammatory markers | 48
open wound | 48
draining purulent fluid | 48
aspiration | 48
Musculoskeletal Infection Society | 48
prosthetic joint infection | 48
biopsy | 48
culture | 48
left thigh mass | 48
necrotic tissue | 48
coagulated blood | 48
foul smell | 48
extensive coagulated blood | 48
necrotic tissue | 48
proximal femur | 48
bone loss | 48
prosthesis | 48
acetabular component | 48
friable bone | 48
cup | 48
tissue | 48
pelvis | 48
biopsy | 48
culture | 48
hemostasis | 48
thrombin spray | 48
argon laser | 48
gel foam sponges | 48
Bovie electrocautery | 48
negative-pressure wound therapy | 48
IR | 48
embolization | 48
profunda femoris | 48
medial femoral circumflex arteries | 48
intensive care unit | 48
intubated | 48
extubated | 48
infectious disease consultation | 48
antibiotic regimen | 48
admitting blood cultures | 48
negative | 48
finalized | 48
tumor board conference | 48
differential diagnosis | 48
chronic infection | 48
particle-associated periprosthetic osteolysis | 48
Gorham vanishing bone disease | 48
lymphangioma | 48
vascular tumor | 48
paraneoplastic abdominal tumor | 48
left hemipelvis | 48
nonreconstructable | 48
left hip disarticulation | 48
antibiotics | 48
sitting function | 48
left hemipelvectomy | 48
acetabular component | 96
grossly loose | 96
blunt dissection | 96
serosa | 96
cup | 96
rongeurs | 96
curettes | 96
necrotic tissue | 96
gluteus maximus | 96
polydioxanone suture | 96
drain | 96
anterior | 96
posterior | 96
skin | 96
approximated | 96
staple closure | 96
incisional wound vacuum | 96
CT abdomen and pelvis | 96
gastrointestinal malignancy | 96
left inguinal | 96
pelvic sidewall | 96
para-aortic | 96
retroperitoneal lymphadenopathy | 96
IV cefepime | 96
oral Flagyl | 96
postoperative course | 96
routine healing | 96
antibiotic regimen | 96
oral chronic suppression therapy | 96
linezolid | 96
cefpodoxime | 96
draining wound | 672
posterolateral aspect | 672
incision | 672
wet-to-dry dressing changes | 672
oral antibiotic suppression | 672
conservative chronic antibiotic suppression | 672
wound care | 672
colonoscopy | 672
outpatient gastroenterology | 672
lost to follow-up | 1008
emergency room | 1008
continued wound drainage | 1008
hip incision | 1008
imaging | 1008
left against medical advice | 1008
orthopaedics team | 1008