28 years old | 0
female | 0
admitted to the hospital | 0
intermittent fever | -672
systemic rashes | -120
oral ulcer | -120
edema in both eyelids | -120
cough | -120
sticky white phlegm | -120
red rash | -120
no chills | -672
no cough | -672
no expectoration | -672
no fatigue | -672
no night sweating | -672
antibiotic treatment | -672
poor outcome | -672
body temperature 36.8°C | 0
pulse 110 bpm | 0
respiration 18 bpm | 0
blood pressure 107/79 mmHg | 0
oxygen saturation 97% | 0
conscious but slow responses | 0
limited speech | 0
red rash on face, neck, and limbs | 0
dermohemia on hands and feet | 0
swollen eyelids | 0
weak breathing sounds in lower lungs | 0
heart rate 110 bpm | 0
no tenderness in abdomen | 0
no sifting dullness | 0
no joint tenderness | 0
no neck rigidity | 0
pitting edema in four extremities | 0
WBC count 1.4 × 10^9/L | 0
hemoglobin 89.9 g/L | 0
PLT count 88.5 × 10^9/L | 0
blood in urine 3+ | 0
urine protein 3+ | 0
erythrocyte sedimentation rate 70 mm/hour | 0
C-reactive protein 3.06 mg/L | 0
blood urea nitrogen 12.4 mmol/L | 0
serum creatinine 124.6 µmol/L | 0
serum albumin 20.9 g/L | 0
immunoglobulin A 1.34 g/L | 0
immunoglobulin G 19.10 g/L | 0
immunoglobulin M 1.29 g/L | 0
compliment C3 0.18 g/L | 0
compliment C4 0.13 g/L | 0
antinuclear antibody (+) 1:1280 | 0
anti-ds-DNA antibody (+) 1:160 | 0
anti-histone antibody 183.64 RU/mL | 0
anti-nucleosome antibody 339.34 RU/mL | 0
perinuclear anti-neutrophil cytoplasmic antibodies (+) 1:40 | 0
extractable nuclear antigen antibodies (+) | 0
anti-Smith antibody (+) | 0
methylprednisolone 80 mg twice a day | 0
meropenem | 0
r-globulin 20 g/day | 0
temperature returned to normal | 24
rash faded | 24
cough persisted | 24
expectoration persisted | 24
WBC count increased | 24
PLT count increased | 24
systemic convulsions | 144
loss of consciousness | 144
cyanosis | 144
upturned eyes | 144
trismus | 144
foaming at the mouth | 144
urinary incontinence | 144
sedation | 144
antiepileptic medication | 144
corticosteroids | 144
fever | 144
rapid heart rate | 144
seizure recurred | 168
transferred to intensive care unit | 168
corticosteroids | 168
antiepileptic medication | 168
antipyretic medication | 168
acid suppression medication | 168
electrolyte disorder correction | 168
regained consciousness | 240
loss of consciousness | 288
MRI of head | 288
abnormal signal with shadows in bilateral frontal, parietal, temporal, and occipital lobes | 288
cerebrospinal fluid with elevated protein levels | 288
epilepsy | 288
posterior cerebral encephalopathy syndrome | 288
methylprednisolone 1000 mg once a day | 288
dexamethasone | 288
prednisone tablets | 288
hydroxychloroquine sulfate | 288
cyclophosphamide | 288
r-globulin | 288
symptomatic and supportive therapies | 288
regained consciousness | 312
condition improved | 312
discharged from hospital | 432
MRI of head | 744
lesions mostly absorbed | 744
prednisone tablets 5 mg orally | 744
hydroxychloroquine 0.3 g once a day | 744
mycophenolate mofetil 0.75 g once a day | 744
stable condition | 744