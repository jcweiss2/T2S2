80 years old | 0
woman | 0
admitted to the hospital | 0
abdominal pain | 0
vomiting |#0x0a
