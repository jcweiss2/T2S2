44 years old | 0
male | 0
bronchobiliary fistula | 0
pneumonia | 0
pancreaticoduodenectomy (Whipple operation) | -2928
transarterial embolization | -2928
pseudoaneurysm rupture of the gastroduodenal artery | -2928
dilation of the bile duct | -720
small-sized multiple bilomas in hepatic segment VIII | -720
poor oral intake | -720
fluctuating fever | -720
jaundice | -720
intravenous antibiotic treatment | -720
repeated drainage endoscopic (ERBD) | -720
percutaneous (PTBD) drainage | -720
recurrent biliary stent obstruction | -168
acute dyspnea | -168
yellowish sputum | -168
sputum positive for bilirubin | -168
preoperative chest X-ray | 0
progressive consolidation | 0
pleural effusion in the right lung | 0
abdominal computed tomography (CT) | 0
dilated bile duct | 0
bilomas of various sizes in liver | 0
chest CT | 0
subdiaphragmatic abscess | 0
pneumonic consolidation with necrotizing change in the right lower lung | 0
bilateral pleural effusion | 0
tubogram | 0
fistulous communication between the dilated intrahepatic bile duct and right lower lung | 0
fiberoptic bronchoscopy (FOB) | 0
copious bile originated from the right lower bronchus | 0
preoperative arterial blood gas analysis (ABGA) | 0
pH 7.41 | 0
PaCO2 32 mmHg | 0
PaO2 67 mmHg | 0
HCO3- 20.1 mmol/L | 0
leukocytosis (15,300 /mm3) | 0
total bilirubin 3.74 mg/dL | 0
direct bilirubin 2.30 mg/dL | 0
alkaline phosphatase 560 IU/L | 0
γ-glutamyl transferase 128 U/L | 0
albumin 2.8 g/dL | 0
lactate 2.8 mmol/L | 0
international normalized ratio of prothrombin time 1.57 | 0
Staphylococcus aureus | 0
Escherichia coli | 0
Enterococcus faecium | 0
Pseudomonas aeruginosa | 0
gradual deterioration | 0
hypoxemia | 0
uncontrolled pneumonia | 0
PTBD for preoperative biliary decompression | 0
icteric | 0
productive cough | 0
yellowish sputum | 0
no significant dyspnea | 0
semi-Fowler position | 0
electrocardiogram | 0
pulse oximetry | 0
continuous invasive arterial blood pressure (ABP) | 0
oxygen saturation (SpO2) 94% | 0
heart rate 117 beats/min | 0
ABP 121/75 mmHg | 0
preoxygenated with 100% oxygen | 0
rapid sequence induction | 0
etomidate 6 mg | 0
rocuronium 60 mg | 0
left-sided double-lumen endobronchial tube (DLT) | 0
both lungs ventilated with 50% oxygen | 0
propofol | 0
remifentanil | 0
bispectral index range 40 to 60 | 0
central venous pressure (CVP) | 0
esophageal temperature | 0
urine output | 0
bile-stained secretions | 0
secretions minimal in left bronchus | 0
biliary spillage from right lower bronchus | 0
OLV initiated | 0
tidal volume 8 ml/kg | 0
respiratory rate 15/min | 0
100% oxygen | 0
positive end-expiratory pressure 5 cmH2O | 0
lateral decubitus position | 0
SpO2 decreased to 92% | 0
SpO2 increased to 97% | 0
pH 7.25 | 0
PaCO2 47 mmHg | 0
PaO2 92 mmHg | 0
HCO3− 20.6 mmol/L | 0
bronchial lavage | 0
resection of the fistula | 0
bilobectomy of the right lung | 0
multiple abscess pockets | 0
necrotizing pneumonia | 0
perforated diaphragm | 0
subphrenic drain | 0
oxygenation gradually improved | 0
two-lung ventilation (TLV) reinstituted | 0
recruit maneuver | 0
PaO2 201 mmHg | 0
anesthesia duration 445 minutes | 0
operation duration 340 minutes | 0
estimated blood loss 1 L | 0
ABP 100/60 to 125/70 mmHg | 0
CVP 5 to 10 mmHg | 0
crystalloid 4.2 L | 0
packed red blood cells 2 units | 0
dopamine 3 to 5 μg/kg/min | 0
urine output 1480 mL | 0
hypokalemia | 0
intravenous potassium repletion | 0
DLT replaced with single-lumen endotracheal tube | 0
postoperative mechanical ventilation | 0
sedation with dexmedetomidine | 0
postoperative chest X-ray | 0
decreased effusion of right lung | 0
extubated on the 4th postoperative day | 96
no sign of BBF recurrence | 96
succumbed to progressive sepsis | 2904
wound infection | 2904
hepatic failure | 2904
necrotizing pneumonia | 2904
repeated biliary stent stricture | 2904
