40 years old|0
male|0
presented to the accident and emergency department|0
severe diffuse abdominal pain|0
abdominal bloating|0
diarrhea|0
nausea|0
past medical history of two episodes of acute diverticulitis over the past 2 years|0
hospitalized for a ruptured diverticulum in the sigmoid colon| -87600
temperature 38.8°C|0
heart rate 120 beats/min|0
normal blood pressure|0
normal oxygen saturation|0
abdominal distension|0
tenderness on deep palpation on the left lower quadrant|0
absence of peritoneal signs|0
rectal examination revealed no stool in the vault|0
hemoglobin 15.9 g/dl|0
WBC 19.120|0
NEUT 80.2%|0
CRP 270.6 mg/l|0
CPK 543 U/l|0
GLU 125 mg/dl|0
LDH 481 U/l|0
fibrinogen 4.4 g/l|0
Na 141 mEq/l|0
K 5.2 mEq/l|0
abdominal CT scan showed located stenosis of the sigmoid colon|0
marked dilation of the descending colon (12 cm diameter)|0
dilation of the transverse colon (7.5 cm diameter)|0
dilation of the ascending colon (12 cm diameter)|0
dilation of the cecum (11 cm diameter)|0
prior CT scan showed stenotic lesion in the sigmoid colon with mechanical obstruction and prestenotic dilation of the colon| -17520
prior admission due to acute diverticulitis 2 years earlier| -17520
prior admission due to a crisis of acute diverticulitis 2 years earlier| -17520
mild periodic discomfort in the abdomen| -17520
patient deteriorated over 8 h|8
signs of sepsis|8
multiorgan failure|8
severe dyspnea|8
metabolic acidosis|8
CT scan ruled out pulmonary embolism|8
intubated due to respiratory muscle fatigue|8
CRP 318 mg/l|8
CPK 543 U/l|8
fibrinogen 6 g/l|8
creatinine 2.2 mg/dl|8
PT 28.20 s|8
INR 2.56|8
D-dimer 2,223.2 μg/l|8
Na 133 mEq/l|8
K 5.4 mmol/l|8
P 5.4 mg%|8
compatible with toxic megacolon|8
surgical assessment performed|8
emergency laparotomy decided|8
surgery revealed extensive necrotic colon|8
total colectomy implemented|8
protective loop ileostomy|8
transferred to intensive care unit due to hemodynamic instability|8
extubated after 12 h|20
transferred to the ward|20
discharge 10 days later|248
histological examination revealed resolving necrotic colon|0
specimen negative for malignancy|0
loop ileostomy reversed 3 months later|2184
patient remains in good health today, 4 years later|35064
prior episodes of acute diverticulitis over the past 2 years| -17520
ruptured diverticulum in the sigmoid colon 10 years prior| -87600
refusal of surgery| -87600
conservatively treated| -87600
stenotic lesion in the sigmoid colon with mechanical obstruction| -17520
prestenotic dilation of the colon| -17520
mild periodic discomfort in the abdomen before latest admission| -17520
severe abdominal pain started 8 h earlier| -8
deterioration over 8 h|8
no stool in the vault|0
no pulmonary embolism|8
respiratory muscle fatigue|8
hemodynamic instability|8
discharge after 10 days|248
ileostomy reversal after 3 months|2184
good health 4 years later|35064
