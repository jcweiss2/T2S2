20 years old | 0 | 0 
male | 0 | 0 
non-smoker | 0 | 0 
occupational smoke exposure | -336 | 0 
fever | -336 | 0 
productive cough | -336 | 0 
night sweats | -336 | 0 
malaise | -336 | 0 
myalgia | -336 | 0 
treated with roxithromycin | -168 | -24 
temperature 38.4°C | 0 | 0 
blood pressure 130/70 mmHg | 0 | 0 
pulse 88 bpm | 0 | 0 
oxygen saturation 97% | 0 | 0 
dyspnoea | 0 | 0 
tachypnoea | 0 | 0 
bronchial breathing sounds | 0 | 0 
crackles over the right lung | 0 | 0 
white blood cells 11.54×10^3/μl | 0 | 0 
total eosinophils 92×10^4/μl | 0 | 0 
haemoglobin 13.7 g/dl | 0 | 0 
creatinine 1.1 mg/dl | 0 | 0 
C-reactive protein (CRP) 11 mg/dl | 0 | 0 
liver enzymes elevated | 0 | 0 
ALP 524 | 0 | 0 
GGT 320 | 0 | 0 
ALT 406 | 0 | 0 
AST 137 | 0 | 0 
abdominal ultrasound normal | 0 | 0 
infiltrates involving most of the right lung | 0 | 0 
treated with IV cefuroxime | 0 | 48 
blood and sputum cultures negative | 0 | 48 
urine Legionella antigen test negative | 0 | 48 
high-grade fever | 48 | 96 
antibiotic treatment changed to moxifloxacin | 48 | 48 
respiratory distress | 96 | 120 
oxygen saturation dropped to 88% | 96 | 96 
arterial blood gas disclosed PaO2 67 mmHg | 96 | 96 
CRP increased to 14 mg/dl | 96 | 96 
liver enzymes elevated | 96 | 96 
leucocytosis 12.8×10^3/μl | 96 | 96 
eosinophil count 1.33×10^3 cells/μl | 96 | 96 
diffuse bilateral infiltrates | 96 | 96 
respiratory distress worsened | 120 | 120 
intubated | 120 | 120 
mechanically ventilated | 120 | 120 
transferred to the intensive care unit | 120 | 120 
broncho-alveolar lavage demonstrated 30% eosinophils | 144 | 144 
diagnosis of AEP | 144 | 144 
IV glucocorticoids administered | 144 | 144 
prompt improvement | 144 | 168 
resolution of fever | 144 | 168 
successful extubation | 168 | 168 
chest radiogram revealed considerable regression of the bilateral infiltrates | 168 | 168 
eosinophil count dropped to 260 cells/μl | 168 | 168 
discharged | 192 | 192 
oral prednisone 60 mg/day | 192 | 432 
tapering over 3 months | 192 | 432