48 years old | 0
male | 0
hypertension | 0
hyperlipidemia | 0
chronic back pain | 0
lisinopril | 0
atorvastatin | 0
over-the-counter analgesics | 0
central chest pain | 0
feeling of warmth | 0
temperature of 36.4 Celsius | 0
heart rate of 87/minute | 0
blood pressure of 126/73 mm Hg | 0
respiratory rate of 22/minute | 0
oxygen saturation 95% | 0
white blood cell count 9000/cumm | 0
neutrophil count 76.6% | 0
lymphocyte count 15.4% | 0
absolute lymphocyte count 1.40 K/mm | 0
lactic acid level 1.3 mmol/L | 0
erythrocyte sedimentation rate 62 mm/hr | 0
c-reactive protein 8.66 mg/dl | 0
troponin <0.03 ng/ml | 0
procalcitonin 0.19 ng/ml | 0
normal sinus rhythm | 0
no ST changes | 0
no T wave changes | 0
chest x-ray hypo inflation | 0
chest x-ray perihilar air space opacities | 0
chest x-ray atelectasis | 0
bilateral ground glass opacities | 0
blood cultures | 0
sputum culture | 0
viral respiratory panel | 0
ceftriaxone | 0
azithromycin | 0
pneumonia | 0
admitted to general medical floors | 0
tachycardic | -48
hypoxic | -48
continued fevers | -48
tested positive for SARS CoV-2 | -48
evaluated by infectious disease consultant | -48
hydroxychloroquine | -48
non-invasive ventilation | -72
endotracheal intubation | -120
transfer to intensive care unit | -120
ARDS | -120
prone position for 16 hours a day | -120
ST elevations in leads II, III, and aVF | -192
troponin peak 0.10 ng/ml | -192
clopidogrel 300 mg | -192
clopidogrel 75 mg daily | -192
evaluated by Cardiology | -192
acute coronary syndrome | -192
serial ECGs | -216
ST changes resolved | -216
coronary catheterization deferred | -216
focal pericarditis | -216
echocardiogram deferred | -216
intermittent fevers | -192
elevated ESR 122 mm/hr | -192
elevated CRP 17.86 mg/dl | -192
cytokine storm | -192
methylprednisolone 1 mg/kg | -192
dexamethasone 20 mg daily | -192
dexamethasone tapered off over 21 days | -192
convalescent plasma candidate | -192
deep vein thrombosis | -216
prophylactic anticoagulation | -216
therapeutic anticoagulation | -216
intravenous plasma | -216
critical respiratory status | -216
echocardiogram normal left ventricular function | -336
no regional wall motion abnormalities | -336
inpatient | 0
discharged | N/A
