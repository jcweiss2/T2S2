42 years old | 0\
female | 0\
granular dystrophy | 0\
DALK | 0\
big bubble technique | 0\
infiltrates along the graft-host junction | 24\
severe anterior chamber reaction | 24\
postoperative keratitis | 24\
graft removed | 24\
stromal graft | 24\
corneal scrapings | 24\
microbiology | 24\
host DM clear | 24\
intact | 24\
residual infiltrates | 24\
topical vancomycin | 27\
topical ceftazidime | 27\
Gram-negative Bacilli | 48\
infiltrates along the entire graft host junction | 48\
hypopyon | 48\
topical antibiotics | 48\
Klebsiella pneumoniae | 48\
resistant to cefazolin | 48\
resistant to amikacin | 48\
resistant to vancomycin | 48\
resistant to ceftazidime | 48\
resistant to ofloxacin | 48\
resistant to ciprofloxacin | 48\
resistant to moxifloxacin | 48\
resistant to cefixime | 48\
resistant to chloramphenicol | 48\
resistant to tetracycline | 48\
resistant to gentamicin | 48\
resistant to cefalexin | 48\
sensitive to imipenem | 48\
sensitive to tigecycline | 48\
partially sensitive to gatifloxacin | 48\
imipenem drops | 48\
infiltration extended | 72\
hypopyon persisted | 72\
therapeutic penetrating keratoplasty | 96\
infiltrates in host DM | 96\
graft clear | 120\
infiltrates resolved | 120\
hypopyon resolved | 120\
gatifloxacin drops | 120\
prednisolone drops | 144\
unaided vision 6/60 | 432\
pin hole vision 6/18 | 432\
graft clear | 432\
anterior segment quiet | 432\
intraocular pressure normal | 432\
pathogen eradicated | 432