56 years old | 0
male | 0
diarrhea | -480
yellow loose stools | -480
diarrhea aggravated | -240
dark green watery stool | -240
palpitations | -240
shortness of breath | -240
dizziness | -240
dry mouth | -240
dry skin | -240
sunken eye socket | -240
no fever | -168
no abdominal pain | -168
no traveling | -168
allograft | -17544
tacrolimus | -17544
mycophenolic acid | -17544
sirolimus | -17544
temperature 37.9°C | 0
septic shock | 0
metabolic acidosis | 0
intubated | 0
transferred to ICU | 0
oliguria | 0
serum creatinine 170 μmol/L | 0
acute kidney injury | 0
CRRT | 0
WBC count 13.46×10^9/L | 0
elevated neutrophil ratio 87.9% | 0
PCT 3.32 ng/mL | 0
CRP 190 mg/L | 0
TPN-T 191.2 ng/L | 0
no significant changes in liver function | 0
no significant changes in blood coagulation | 0
no significant changes in platelet count | 0
tacrolimus within target range | 0
temperature rise to 38.5°C | 24
piperacillin/tazobactam | 24
bronchoalveolar lavage culture | 24
Aspergillus fumigatus | 24
carbapenem-resistant Klebsiella pneumoniae | 24
urine bacterial culture negative | 24
venous blood culture negative | 24
anaerobic blood culture negative | 24
meropenem | 24
voriconazole | 24
tacrolimus discontinued | 24
sirolimus discontinued | 24
stool detection | 24
intestinal bacterial culture negative | 24
parasite microscopic exam negative | 24
clostridium difficile antigen negative | 24
compound berberine | 24
correct electrolyte balance | 24
correct acid-base balance | 24
diarrhea mitigated | 24
enteral nutrition solution | 24
probiotics | 24
high frequency diarrhea | 48
fever 39°C | 48
parasitic stool exam negative | 48
fecal bacterial culture negative | 48
blood mNGS analysis | 48
Klebsiella pneumoniae | 72
Cryptosporidium parvum | 72
Cryptosporidium oocysts | 72
azithromycin | 72
liver function indices elevated | 72
T lymphocyte count elevated | 72
cyclosporine added | 72
cyclosporine trough 194.00 μg/L | 96
cyclosporine dose adjusted | 96
azithromycin stopped | 168
nitazoxanide added | 168
diarrhea frequency reduced | 216
diarrhea subsided | 336
Cryptosporidium oocysts absent | 336
nitazoxanide stopped | 336
systemic infection controlled | 960
disconnected from ventilator | 960
creatinine normalized | 960
liver function recovered | 960
condition stabilized | 1128
no ventilator reliance | 1128
transferred to general ward | 1128
