48 years old | 0
male | 0
high grade urothelial carcinoma | -40320
carcinoma in situ | -40320
radical cystectomy | -40320
orthotopic Studer ileal neobladder | -40320
right laparoscopic nephroureterectomy | -17520
upper urinary tract urothelial carcinoma | -17520
referred to emergency department | 0
impaired kidney function | 0
serum creatinine 3.5 mg/dL | 0
no flank pain | 0
no gross hematuria | 0
no fever | 0
clean intermittent self-catheterization every 4 hours | 0
denied decreased output of urine | 0
urinary catheter placed | 0
serum creatinine 4 mg/dL | 0
renal ultrasound revealed severe hydronephrosis | 0
computed tomography (CT) scan performed | 0
smooth-walled stricture of distal left ureter | 0
severe dilatation of urinary tract above stricture | 0
empty Studer-type neobladder | 0
presumptive diagnosis benign ureteroileal stricture | 0
10F percutaneous nephrostomy (PN) tube placed | 0
shaking chills | 24
tachycardia | 24
septic shock | 24
anesthesia consulted | 24
hemodynamic support | 24
discharged from intensive care unit (ICU) | 48
multifactorial acute kidney failure | 48
serum creatinine around 8 mg/dL | 48
favourable follow-up after ICU discharge | 48
episode of massive and life-threatening hematuria | 168
important bleeding through PN tube (approximately 700ml) | 168
urgent CT angiography performed | 168
renal pseudoaneurysm of segmental renal artery | 168
hyperdense material indicative of blood clots in collecting system | 168
superselective endovascular embolization with Onyx® performed | 168
exclusion of pseudoaneurysm | 168
prior hemoglobin level 12.8 g/dL | 168
hemoglobin dropped to 7.2 g/dL | 168
transfusion of 2 RBC units | 168
hemoglobin increased to 9 g/dL | 168
hemoglobin stable at discharge | 168
urine remained clear | 168
renal function progressively improved | 168
serum creatinine 3 mg/dL | 168
