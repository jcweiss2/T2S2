30 years old | 0
G1P0 | 0
Hispanic female | 0
presented at 15 weeks gestation | 0
acute right lower quadrant abdominal pain | -120
acute right upper quadrant abdominal pain | -120
progressive right lower quadrant abdominal pain | -120
progressive right upper quadrant abdominal pain | -120
dysuria | -120
nausea | -120
vomiting | -120
emesis progressed to complete oral intolerance | -132
emergency department presentation 3 days prior | -168
acute hyperemesis gravidarum | -168
obstetrical ultrasound | -168
single living intrauterine pregnancy | -168
estimated gestation age of 13 weeks | -168
fetal heart tones measured 160 bpm | -168
no mention of appendiceal imaging | -168
orally challenged successfully | -168
discharged home with oral antibiotics | -168
discharged home with antiemetics | -168
abdominal pain in the right lower quadrant | 0
abdominal pain in the right upper quadrant | 0
abdominal pain in the left lower quadrant | 0
moderate tenderness to palpation in the right lower quadrant | 0
white blood cell count increased to 16200 | 0
ultrasound imaging revealed dilated fluid filled bowel | 0
fetal heart tones reported at 160 bpm | 0
acute gestational appendicitis diagnosed | 0
general surgery consultation requested | 0
clinical diagnosis confirmed | 0
laparoscopic abdominal access achieved | 0
massive bowel distention | 0
purulent ascites | 0
conversion from laparoscopy to open laparotomy | 0
abscess discovered enveloping the ileocecum | 0
perforation of the appendiceal base | 0
extension into the cecum | 0
cecal necrosis | 0
ileocecectomy performed | 0
abdomen irrigated | 0
attempted fascial closure abandoned | 0
significant abdominal wall tension | 0
pronounced bowel edema | 0
ACS diagnosed | 0
abdomen left open | 0
temporary closure performed using sterile radiologic cassette cover | 0
perforated with #10 blade scapel | 0
saline-dampened surgical towel placed | 0
two 10-French flat surgical drains | 0
closure of the abdominal domain with loban drape | 0
intubated | 0
transferred to ICU | 0
intravenous antibiotics | 0
resuscitation fluids | 0
consultations with infectious disease | 0
consultations with obstetrician | 0
daily fetal heart tones determined | 0
negative pressure therapy maintained at 120–130 mmHg | 0
peritoneal toilet performed on post-operative day 4 | 96
inspection of the ileocolic anastomosis | 96
complete integrity | 96
no evidence of bowel necrosis | 96
significant bowel edema | 96
temporary abdominal closure achieved | 96
fascial closure achieved on post-operative day 6 | 144
skin closure deferred | 144
wound VAC with GRANUFOAM | 144
extubated in ICU | 144
delayed primary closure of laparotomy incision on post-operative day 12 | 288
progressed to regular diet | 288
pathology diagnosis of acute ruptured appendicitis | 288
abscess formation | 288
acute serositis | 288
discharged home on post-operative day 15 | 360
tocolysis not indicated | 360
deferred throughout admission | 360
eventual normal spontaneous vaginal delivery | 0
no incisional hernia development at 5 years | 0
daughter obtained all developmental milestones | 0
developed only common childhood illnesses | 0
