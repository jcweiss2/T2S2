27 years old | 0
female | 0
Caucasian | 0
admitted to the hospital | 0
history of intravenous drug use | -2160
tricuspid valve endocarditis | -2160
bacteraemia | -2160
Candida | -2160
Staphylococcus aureus | -2160
treated with 6 weeks of IV antibiotics | -2160
treated with anti-fungals | -2160
vancomycin | -2160
daptomycin | -2160
linezolid | -2160
cefepime | -2160
micafungin | -2160
tricuspid valve replaced with CorMatrix extracellular-based material | -2160
post-operative complications of pulmonary embolism | -2160
Coumadin initiated | -2160
surveillance blood cultures returning positive for methicillin-sensitive S. aureus | 0
surveillance blood cultures returning positive for Candida parapsilosis | 0
gingival haemorrhage | 0
spontaneous bruising | 0
abdominal swelling | 0
supratherapeutic international normalized ratio | 0
thrombocytopenia | 0
computed tomography abdomen and pelvis showed large pericardial effusion | 0
hepatosplenomegaly | 0
mild ascites | 0
infectious disease consulted | 0
nafcillin initiated | 0
amphotericin B initiated | 0
admitted to the Cardiology Intermediate Unit | 0
echocardiogram shows large mobile mass involving the TV | 24
echocardiogram shows large pericardial effusion | 24
evidence of markedly elevated intrapericardial pressure | 24
causing diastolic compression of the right ventricle | 24
ultrasound-guided pericardiocentesis | 24
removal of 600 mL of serous fluid | 24
echocardiogram showed residual moderate effusion | 48
nafcillin switched to cefazolin | 48
amphotericin B continued | 48
blood cultures from 02/13 return positive for Mycobacteria | 72
amphotericin B discontinued | 72
switched to fluconazole | 72
echocardiogram shows severe TV thickening | 72
large vegetation is pedunculated and mobile | 72
ruptured TV chordae | 72
flail septal leaflet | 72
effusion measures 2.8 cm anteriorly and 3.8cm posteriorly | 72
evidence of right ventricular compression | 72
blood cultures from 02/18 return positive for C. parapsilosis | 168
clinical deterioration | 168
tachycardia | 168
increased dyspnoea | 168
abdominal distension | 168
lower extremity oedema | 168
persistent fevers | 168
lactic acid at nine | 168
transferred to the CICU | 168
echocardiogram shows severe ‘torrential’ wide open tricuspid regurgitation | 168
flail septal leaflet of TV | 168
echodensity attached to tip suggestive of ruptured chordae and/or vegetation | 168
large vegetation attached to tricuspid leaflet is no longer visualized | 168
suspicious for embolization | 168
cefazolin and fluconazole switched to liposomal amphotericin B | 168
amikacin initiated | 168
imipenem initiated | 168
azithromycin initiated | 168
continued clinical deterioration | 192
tachypneic | 192
hypoxic | 192
hypotensive | 192
requiring intubation | 192
requiring pressors | 192
continued clinical decline | 216
severe metabolic acidosis | 216
lactic acid of 19 | 216
pH of 7.27 | 216
signs of multiorgan failure | 216
taken to the OR for emergent TVR | 216
emergency redo sternotomy | 216
redo TV replacement with 29 Biocor valve | 216
removal of embolized old CorMatrix TV from right pulmonary artery | 216
blood cultures from 02/19 return positive for Mycobacterium | 240
amphotericin B switched to micafungin | 240
amikacin continued | 240
imipenem continued | 240
azithromycin continued | 240
recommendations to complete micafungin for a total of 6 weeks | 240
recommendations to complete antibiotics for a total of 3 months | 240
patient discharged home | 672
Linezolid initiated | 672
Amikacin initiated | 672
Micafungin initiated | 672
all laboratory values improved | 672
patient moved out of state | 672
re-admitted within 2 months | 1344
blood cultures positive for AFB | 1344
TEE revealed new TV vegetations | 1344
recurrent IVDU | 1344
not a candidate for surgical intervention | 1344
treated with 6 weeks of Linezolid | 1344
treated with Imipenem | 1344
lost to follow-up | 1344