69 years old | 0
man | 0
history of ischaemic heart disease | 0
history of chronic liver disease | 0
history of adrenal incidentaloma | 0
history of arterial hypertension | 0
history of diabetes mellitus type 2 | 0
history of hyperuricaemia | 0
history of dyslipidaemia | 0
hospital admissions (four in previous 5 months) | -3600
bacteraemia caused by ESBL-producing Escherichia coli | -3600
bacteraemia caused by Klebsiella pneumoniae | -3600
unknown focus of infection | -3600
fever | 0
dyspnoea | 0
dizziness | 0
diffuse abdominal pain | 0
Murphy’s sign absent | 0
elevated plasma C-reactive protein | 0
elevated plasma procalcitonin | 0
blood culture negative | 0
heterogeneous liver (ultrasound) | 0
cholelithiasis | 0
focus of infection in gallbladder and biliary tract hypothesis | 0
laparoscopic cholecystectomy | 0
hepatic lesions identified | 0
hepatic lesions biopsied | 0
calcified biliary hamartomas (histology) | 0
K. pneumoniae confirmed (bacteriology) | 0
clinical improvement | 24
discharged | 24
re-admitted to intensive care unit | 720
bacteraemia due to ESBL-producing K. pneumoniae | 720
abdominal contrast-enhanced CT scan | 720
liver with increased dimensions | 720
liver heterogeneous texture | 720
multiple calcified lesions (related to granulomas) | 720
hypodense area (24 mm) in left lobe (segment III) | 720
MRI | 720
several nodular lesions | 720
probable calcifications | 720
largest lesion (2.8 cm) | 720
morphological alteration of liver with evident hypertrophy | 720
chronic hepatopathy | 720
hepatobiliary scintigraphy | 720
bile ducts normal appearance | 720
no obstruction | 720
recurrent sepsis | 720
multidisciplinary meeting | 720
liver transplant ruled out | 720
MRI benign lesions | 720
absence of hepatic cirrhosis signs | 720
broad-spectrum antibiotics cycles | 720
meropenem 1g three times a day (14 days) | 720
amikacin 500mg twice a day (17 days) | 720
piperacillin and tazobactam 4.5g four times a day (17 days) | 720
ceftriaxone 1g once a day (10 days) | 720
favourable clinical evolution | 720
improvement after each cycle | 720
discharged at treatment completion | 720
readmitted again (four months after surgery) | 2880
sepsis | 2880
bacteraemia due to ESBL-producing K. pneumoniae | 2880
focus of infection hypothesized as biliary hamartomas | 2880
extended cycle of meropenem 1g three times a day (21 days) | 2880
discharged after 3 weeks | 2880
prophylactic antibiotics | 2880
surveillance by consultant | 2880
no relapse (3 years follow-up) | 26280
no symptoms related to previous admissions | 26280
prophylactic antibiotic (ciprofloxacin 500mg twice a day) | 26280
annual MRI | 26280
