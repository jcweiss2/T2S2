68 years old| 0
    female | 0
    admitted to the hospital | 0
    AML | -4320
    bone marrow biopsy (80% blasts) | -4320
    white blood cell count 175,000 | -4320
    27% peripheral blasts | -4320
    normal karyotype on cytogenetics | -4320
    DNMT3 mutation | -4320
    NPM1 mutation | -4320
    PTPN11 mutation | -4320
    TET2 mutations | -4320
    induction chemotherapy (decitabine and venetoclax) | -4320
    nonsustained ventricular tachycardia | -4320
    rapid atrial fibrillation | -4320
    bacterial pneumonia | -4320
    remission | -4320
    maculopapular rash (torso and upper extremities) | -4320
    leukemia cutis | -4320
    44% monocytic blasts | -4320
    nonproductive cough | -4320
    rhinorrhea | -4320
    sore throat | -4320
    afebrile | -4320
    SARS-CoV-2 positive | -4320
    COVID-19 diagnosis | -4320
    mRNA-1273 vaccine (two doses) | -4320
    admitted to medicine service | 0
    computed tomography chest (no pneumonia) | 0
    no supplemental oxygen | 0
    no intubation | 0
    remdesivir (3-day course) | 0
    hemodynamically stable | 0
    resolved upper respiratory symptoms | 0
    SARS-CoV-2 positive | 72
    transferred to malignant hematology service | 72
    7+3 reinduction chemotherapy (cytarabine and idarubicin) | 72
    intrathecal cytarabine (prophylactic) | 72
    retested every 3–5 days for COVID-19 | 72
    sotrovimab | 168
    SARS-CoV-2 positive | 168
    chest pain | 168
    computed tomography chest (pericarditis) | 168
    pericardial effusion | 168
    colchicine (3-month course) | 168
    resolution of chest pain | 168
    blood cell counts nadir (day 9) | 216
    absolute neutrophil count 0 | 216
    neutropenic fever | 480
    asymptomatic | 480
    negative chest x-ray | 480
    cefepime (7-day course) | 480
    valacyclovir prophylaxis | 480
    isavuconazole prophylaxis | 480
    levofloxacin prophylaxis | 480
    counts recovery (ANC 170) | 600
    ANC 170 | 600
    COVID-19 PCR monitoring | 600
    discharge | 864
    bone marrow biopsy (complete remission) | 864
    persistent DNMT3 mutation | 864
    persistent TET2 mutation | 864
    leukemia cutis rash cleared | 864
    COVID-19 PCR negative | 1008
    high-dose cytarabine consolidation | 1008
    tixagevimab/cilgavimab prophylaxis | 1008
    remained SARS-CoV-2 negative | 1008
    no comorbidities | 0
    vaccination | -4320
    resolved COVID-19 symptoms | 72
    no COVID-19 progression during neutropenia | 480
    neutropenic fever (no respiratory symptoms) | 480
    ANC recovery | 600
    viral load decrease | 600
    neutrophil recovery | 864
    cleared SARS-CoV-2 | 1008
    no repeat infection | 1008
    complete morphologic remission | 864
    clearance of mutations | 864
    mild COVID-19 | 0
    immunocompromise | 0
    antiviral treatment | 0
    frequent viral testing | 0
    no progression to propagating phase | 0
    no progression to complicated phase | 0
    NAAT positive | 0
    no septic shock | 0
    no multiorgan failure | 0
    isolation techniques | 0
    personal protective equipment | 0
    no replicating virus | 1008
    AML therapy complications | 72
    no intensive care needed | 72
    excellent performance status | 864
    energy excellent | 864
    leukemia treatment response | 864
    COVID9-19 recommendations | 0
    delay therapy if possible | 0
    lifesaving chemotherapy considered | 0
    mild infection | 0
    medically stable | 0
    vaccinated | -4320
    antiviral monitoring | 0