42 years old | 0
male | 0
admitted to the hospital | 0
upper abdomen paroxysmal cramp | -168
multiple kidney stones | -8760
treated for kidney stones | -8760
excreted a large amount of tarry stool | 48
coffee-ground emesis | 48
blood pressure dropped | 48
received a blood transfusion | 48
rehydration | 48
transferred to the Intensive Care Unit | 48
bedside upper gastrointestinal endoscopy | 48
duodenal ulcer with an adherent clot | 48
intragastric local instillation of norepinephrine | 48
intragastric local instillation of epinephrine | 48
excreted a large amount of tarry stools | 56
vomited a copious amount of coffee-ground material | 56
subtotal gastrectomy | 56
Billroth II gastrointestinal anastomosis | 56
heart rate became rapid | 96
central venous pressure dropped | 96
blood hemoglobin decreased | 96
abdominal circumference increased | 96
ultrasound examination detected a hematocele | 96
gastroduodenal artery embolization | 96
elevated serum calcium level | 96
low serum phosphorus level | 96
renal dysfunction | 96
elevated plasma parathyroid hormone level | 96
neck computed tomography scan | 96
two enhancing masses in the rear of the right lobe of thyroid gland | 96
severe abdominal pain | 120
tenderness | 120
guarding | 120
rebound pain upon abdominal palpation | 120
rapid heart rate | 120
high leucocyte count in blood | 120
peritonitis | 120
sepsis | 120
intravenous antibiotics | 120
imipenem | 120
tigecycline | 120
continuous renal replacement therapy | 120
elective surgical exploration | 456
excision of the parathyroid adenoma | 456
histology of parathyroid gland revealed a typical parathyroid adenoma | 456
normalized PTH level | 528
decreased calcium level | 528
transferred to the general ward | 528
follow-up | 744
denied any digestive tract symptoms | 744