24 years old | 0
    primiparous | 0
    Japanese | 0
    woman | 0
    no significant medical history | 0
    no complications during pregnancy | 0
    gave birth via vaginal delivery | 0
    healthy baby girl | 0
    depressive mood | -504
    emotional incontinence | -504
    auditory hallucination | -408
    abnormal behavior | -408
    mandatorily hospitalized | -408
    postpartum psychosis | -408
    antipsychotic drugs | -408
    somnolence | -384
    unstable breathing | -384
    generalized seizure | -384
    status epilepticus | -360
    hyperthermia | -360
    transferred to ICU | -360
    generalized seizure difficult to control | -360
    respiratory depression | -360
    tracheal intubation | -360
    artificial ventilation | -360
    methylprednisolone pulse therapy | -360
    IVIg therapy | -360
    symptoms deteriorated | -336
    involuntary movements | -336
    transferred to Shinshu University Hospital | -240
    body temperature 38.5°C | 0
    orofacial dyskinesia | 0
    athetoid movement in right hand | 0
    no nuchal stiffness | 0
    no pathological reflexes | 0
    inflammatory reaction | 0
    mild liver dysfunction | 0
    tests negative for herpes simplex | 0
    tests negative for herpes zoster | 0
    tests negative for Epstein-Barr virus | 0
    anti-thyroglobulin antibody positive | 0
    anti-thyroperoxidase antibody positive | 0
    CSF lymphocytic pleocytosis | 0
    CSF slightly elevated protein | 0
    CSF normal glucose | 0
    anti-NMDAR antibody positive | 0
    EEG extreme delta brush | 0
    brain MRI increased signal | 0
    right ovarian cystic tumor | 0
    anti-NMDAR encephalitis diagnosis | 0
    laparoscopic removal of ovarian tumor | 1344
    mature cystic teratoma | 1344
    IVIg | 1344
    mPSL pulse therapy | 1344
    plasma exchange | 1344
    DFPP | 1344
    involuntary movements prolonged | 1344
    higher brain dysfunction prolonged | 1344
    autonomic dysfunction prolonged | 1344
    repetitive severe infections | 1344
    pneumonia | 1344
    sepsis | 1344
    anti-NMDAR antibody decreased | 1344
    involuntary movements improved | 1344
    respiratory failure improved | 1344
    transferred to rehabilitation hospital | 1344
    bedridden state | 1344
    severe cognitive dysfunction | 1344
    brain MRI almost normal | 1344
    neurological condition continued to improve | 1344
    independent gait | 1344
    verbal communication | 1344
    memory disturbance | 1344
    mental juvenility | 1344
    no brain atrophy | 1344
    no abnormal signals | 1344
    <|eot_id|>
    