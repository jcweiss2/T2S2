70 years old | 0
male | 0
non-hypertensive | 0
non-smoker | 0
well-controlled diabetic | 0
HbA1c = 6.83% | 0
admitted to the hospital | 0
unresolving back pain | -144
COVID-19-induced pneumonia | -144
elevated white blood cell count | 0
WBC = 15,200/mm3 | 0
no abnormal monoclonal gammopathy | 0
contrast-enhanced chest-abdomen-pelvis CT | 0
mediastinal calcified lymph nodes | 0
dense infiltrative retroesophageal prevertebral lesion | 0
lung fields clear | 0
retractile subpleural fibrous bands | 0
stepwise increase in WBC | 0
stepwise increase in CRP | 0
broad spectrum antibiotherapy initiated | 0
dorsal MR | 72
expanding prevertebral lesion | 72
Tuberculosis testing negative | 72
HIV testing negative | 72
brucellosis testing negative | 72
blood culture negative | 72
serum galactomannan assay negative | 72
RT-PCR COVID-19 negative | 72
first percutaneous CT-guided biopsy | 72
biopsy inconclusive | 72
rising WBC count | 240
rising CRP | 240
control dorsal MR | 240
slight progression of the lesion | 240
empirical antifungal therapy initiated | 288
fluconazole 400 mg b.i.d. | 288
amphotericin B 400 mg q.d. | 288
second CT-guided biopsy | 290
necrotic lesions containing fungal organisms | 290
acute-angle-branching hyphae | 290
Aspergillus fumigatus culture positive | 290
antifungal therapy switched to voriconazole | 290
voriconazole 400 mg b.i.d. | 290
voriconazole dosage reduced to 200 mg b.i.d. | 294
surgical thoracotomy not executed | 294
CRP levels decreased | 304
increasing levels of creatinine | 304
progressive oliguria | 304
hemodialysis sessions | 304
paraplegia | 360
altered mental state | 360
ICU transfer | 360
head CT | 360
no focal abnormality in brain parenchyma | 360
lumbar puncture normal | 360
sterile cultures | 360
dorsal MR | 360
spinal cord compression | 360
recent spinal cord compression at T6 to T8 | 360
high signal abnormality on T2-weighted images | 360
prevertebral lesion thickness increased | 360
renal function deteriorating | 432
neurological function deteriorating | 432
comatose | 432
intubated | 432
passed away | 504