57 years old | 0
    man | 0
    presented | 0
    generalized weakness | -336
    fatigue | -336
    confusion | -336
    dizziness | -336
    mild jaundice | -336
    hypertension | 0
    diabetes mellitus | 0
    hyperlipidemia | 0
    hypothyroidism | 0
    former smoker | 0
    consumed alcohol occasionally | 0
    anemia | 0
    thrombocytopenia | 0
    acute liver injury | 0
    acute renal failure | 0
    intermittent hemodialysis | 0
    transferred to medical ICU | 0
    lactic acidosis | 0
    sepsis | 0
    worsening hepatic encephalopathy | 0
    febrile | 0
    hemoglobin 7.5 g/dL | 0
    platelets 26,000/mm³ | 0
    creatinine 4.34 mg/dL | 0
    total bilirubin 19 mg/dL | 0
    alanine aminotransferase 395 U/L | 0
    aspartate aminotransferase 261 U/L | 0
    serum lactate 10 mmol/L | 0
    serum ferritin >40,000 ng/mL | 0
    serum triglycerides 556 mg/dL | 0
    coagulopathic | 0
    international normalized ratio 4.2 | 0
    fibrinogen <70 mg/dL | 0
    MELD score >40 | 0
    emergent liver transplant evaluation | 0
    workup for liver failure unrevealing | 0
    computed tomography of abdomen and pelvis | 0
    hepatic steatosis | 0
    no focal hepatic lesions | 0
    splenomegaly | 0
    multiple splenic infarcts | 0
    right axillary lymphadenopathy | 0
    retropectal lymphadenopathy | 0
    mechanical ventilation | 0
    circulatory shock | 0
    vasopressor support | 0
    worsening renal failure | 0
    continuous renal replacement therapy | 0
    bone marrow biopsy | 0
    no evidence of leukemia | 0
    no evidence of lymphoma | 0
    no evidence of HLH | 0
    removed from transplant list | 0
    transjugular liver biopsy | 0
    diffuse large B-cell lymphoma | 0
    met criteria for HLH | 0
    fever | 0
    bicytopenia | 0
    splenomegaly | 0
    ferritin level | 0
    hypertriglyceridemia | 0
    started on chemotherapy | 0
    dexamethasone | 0
    ifosfamide | 0
    carboplatin | 0
    etoposide | 0
    worsening metabolic acidosis | 0
    hypoglycemia | 0
    shock | 0
    subdural hemorrhages | 0
    generalized tonic-clonic seizures | 0
    family decided on comfort care | 0
    died | 120
    

    
    