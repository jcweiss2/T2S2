60 years old | 0
male | 0
admitted to the emergency room | 0
severe epigastric dilation | 0
stomachache | 0
fever | 0
localized epigastric pain | -48
vomiting | -12
abdominal pain spread to entire stomach | -12
high fever of 39.5°C | -12
endoscopic biliary stenting operation | -336
obstructive jaundice | -336
unresectable pancreatic cancer | -336
serum total bilirubin decreased | -336
direct bilirubin decreased | -336
discharge after stenting | -336
blood pressure 95/65 mmHg | 0
pulse 110 bpm | 0
abdominal distention | 0
hepatomegaly | 0
liver span 2 cm below right costal margin | 0
epigastric tenderness | 0
mild rebounding pain | 0
almost no gurgling sound | 0
emergency abdominal CT scan | 0
irregular gas-containing lesions in liver | 0
liver parenchymal moth-eaten destruction | 0
pneumatized bile duct | 0
no obvious inflammation | 0
stent in common bile duct without obstruction | 0
intrahepatic duct dilation due to obstruction of pancreatic mass | 0
severe intrahepatic infection caused by enterogenous aerogenes | 0
multiorgan deficiency | 0
hepatic injury | 0
renal injury | 0
cardiac injury | 0
coagulopathy | 0
board-spectrum antibiotic treatment | 0
biapenem 0.3 g Q12H | 0
ornidazole 100 mg Q12H | 0
vigorous fluid resuscitation | 0
intensive care | 0
blood pressure falling | 10
inotropic support | 10
norepinephrine infusion | 10
clinical condition deteriorated | 10
multiorgan failure | 10
sudden cardiac arrest | 20
death | 20
blood specimen culture | 24
Clostridium perfringens infection confirmed | 24
Clostridium perfringens bacteremia | 24
Clostridium perfringens liver abscess | 24
phospholipase C lecithinase (α-toxin) | 24
β-toxin | 24
ε-toxin | 24
gas gangrene | 24
capillary leakage | 24
advanced pancreatic cancer | -336
palliative therapy | -336
common bile duct stenting complication | -336
