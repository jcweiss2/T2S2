27 years old | 0
male | 0
residing in Kathmandu | 0
admitted to the clinic | 0
fever | -48
axillary temperature 101.8°F | -48
blood pressure 124/80 mmHg | -48
pulse 86 bpm | -48
denied prior comorbidities | -48
thyroid illness | -48
diabetes mellitus | -48
immunocompromised state | -48
review of systems was normal | -48
dengue non-structural protein 1 (NS1) test sent | -48
dengue NS1 test positive | -48
negative IgG/IgM | -48
haemoglobin 16.7 gm/dl | -48
white blood cell (WBC) 6×10^3/mm^3 | -48
platelet 131×10^3/mm^3 | -48
antipyretics | -48
vomiting | -24
severe headache | -24
myalgia | -24
rash | -24
axillary temperature 100.5°F | -24
blood pressure 130/84 mmHg | -24
pulse 92 bpm | -24
petechiae | -24
hospitalized | 0
treated per guidelines | 0
analgesics | 0
antipyretics | 0
bed rest | 0
fluids | 0
nutritional support | 0
WBC and platelets dropped | 144
sharp chest pain | 144
Electrocardiogram | 144
Troponin-I | 144
ultrasonography (USG) | 240
borderline splenomegaly | 240
minimal left-sided pleural effusion | 240
severe pain in lower limbs | 240
fever peaked at 100.4°F | 240
blood pressure 100/80 mmHg | 240
heart rate 97 bpm | 240
focal tenderness in left buttock | 240
left lumbosacral region | 240
bilateral medial thigh | 240
diagnostic investigations | 240
routine examination of urine and stool | 240
cultures of urine, stool, and blood | 240
Human Immunodeficiency virus | 240
Brucella | 240
Scrub Typhus | 240
Typhoid | 240
Malaria | 240
Leptospirosis | 240
NS1 test for dengue | 240
inflammatory markers | 240
erythrocytic sedimentation rate | 240
C-reactive protein | 240
procalcitonin | 240
Creatinine kinase | 240
troponin level | 240
echocardiography | 240
cannula site looked normal | 240
no history of recent trauma | 240
no intramuscular injections | 240
no recreational drug usage | 240
plain MRI of the Lumbosacral Spine | 312
pyomyositis | 312
Clindamycin | 312
Tazobactam-piperacillin | 312
aspiration | 312
purulent fluid | 312
Gram staining | 312
culture grew Methicillin Sensitive Staphylococcus aureus | 312
antibiotics switched to Cloxacillin | 312
Tazobactam-piperacillin | 312
dual intravenous antibiotics | 312
oral Cloxacillin | 312
repeat USG of the left thigh | 432
collection measuring 7.6×3.5×2.1 cm | 432
aspirated ~30 ml of pus-like fluid | 432
subsequent USG examinations | 432
decreasing amount of fluid collection | 432
discharged on oral antibiotics | 600
USG performed at the end of 6 weeks | 1008
absence of any intramuscular collection | 1008