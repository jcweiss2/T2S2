75 years old | 0
female | 0
admitted to the hospital | 0
epigastric pain | -48
right upper quadrant pain | -48
nausea | -48
no fever | -48
nonspecific digestive difficulties | -672
similar episode | -168
cardiorespiratory examination unremarkable | 0
hemodynamically stable | 0
abdomen tender | 0
guarding in the right upper quadrant | 0
positive Murphy's sign | 0
gallbladder distension | 0
wall thickening | 0
2.5 cm stone in the gallbladder lumen | 0
white blood cell count 8.3 × 10^9/l | 0
C-reactive protein 85 mg/l | 0
serum total bilirubin 17.3 µmol/l | 0
alkaline phosphatase 79 IU/l | 0
aspartate aminotransferase 23 IU/l | 0
alanine aminotransferase 29 IU/l | 0
lipase 32 IU/l | 0
sodium 136 mmol/l | 0
potassium 3.8 mmol/l | 0
blood urea 5.1 mmol/l | 0
creatinine 82 µmol/l | 0
troponin I <0.01 U/l | 0
clinical diagnosis acute cholecystitis | 0
ECG showed sinus rhythm | 0
incomplete right branch block | 0
negative T waves in V1–V3 | 0
no sign of ischemia | 0
intravenous antibiotics | 0
fluids | 0
fever | 24
peripheral blood cultures taken | 24
negative peripheral blood cultures | 24
increased white blood cell count | 24
CRP 434 mg/l | 24
normal urea | 24
normal electrolytes | 24
normal liver function | 24
normal amylase | 24
normal bilirubin | 24
planned surgical cholecystectomy | 24
preoperative ECG | 24
ST segment depression in V3 | 24
elevated troponin I level | 24
creatine kinase level 409 U/l | 24
anticoagulation with high-dose low-molecular-weight heparin | 24
aspirin | 24
β-blockers | 24
angiotensin-converting enzyme inhibitors | 24
admitted to the intensive care unit | 24
troponin level decreased | 36
troponin level decreased again | 44
cardiac ultrasound | 48
mildly enlarged right ventricle | 48
no enlargement of the left ventricle | 48
good ejection fraction | 48
right overload septal motion abnormality | 48
pulmonary hypertension | 48
angio-CT | 48
no pulmonary embolism | 48
coronary angiography | 72
no abnormality | 72
normal left ventricular function | 72
abdominal CT | 72
confirmed cholecystitis | 72
excluded empyema or abscess complications | 72
discharged | 168
elective surgery for symptomatic cholelithiasis | 168