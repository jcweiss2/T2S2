59 years old | 0
    female | 0
    admitted to the hospital | 0
    type-1 diabetes | -175200
    end-stage renal failure | -175200
    combined kidney-pancreas transplant | -175200
    second kidney transplant | -62400
    mycophenolate mofetil | -62400
    tacrolimus | -62400
    immunosuppressive regimen | -62400
    intravenous antibiotics | -240
    no clinical improvement | -240
    normal creatinine level | 0
    glycemia within normal range | 0
    bilateral pleural effusion | 0
    bilateral pneumonia | 0
    multiple abdominal intussusceptions | 0
    discontinued immunosuppressive treatment | 0
    exploratory laparotomy | 0
    free intra-abdominal liquid | 0
    4 sites of intussusception | 0
    intramural lesion | 0
    post-transplant lymphoproliferative disorder suspected | 0
    biopsy | 0
    manual desinvagination | 0
    low-grade tubulovillous adenoma | 288
    new episode of bowel obstruction | 288
    CT scan showing 1 intussusception | 288
    progression of pulmonary infection | 288
    operating room | 288
    recurrence of intussusception | 288
    segmental resection indicated | 288
    hemodynamic instability | 288
    septic shock | 288
    vasoactive support | 288
    manual reduction | 288
    no clinical improvement | 288
    multiple organ failure | 408
    died | 432
    multiple tubulovillous adenomas | 432
    necrosis of pancreas graft | 432
    thrombosis of pancreatic artery | 432
    pulmonary adenocarcinoma | 432
    multiple bilateral pulmonary metastases | 432
    lymphangitic carcinomatosis | 432
    