3 years old | 0
    boy | 0
    admitted | 0
    cough | -48
    cold | -48
    fever | -48
    poor oral intake | -48
    febrile convulsions | -8760
    vomiting | -8760
    cyanosis | -8760
    moderate to high-grade fever | -8760
    deviation of eyes to one side | -8760
    loss of consciousness | -8760
    electroencephalogram (EEG) | -8640
    cerebrospinal fluid studies | -8640
    neuroimaging | -8640
    diagnosis of atypical febrile convulsions | -8640
    no family history of epilepsy | 0
    febrile | 0
    mild congestion in the throat | 0
    symptomatic treatment | 0
    high-grade fever | 4
    vomiting | 4
    bluish discoloration of the extremities | 4
    tachypnea | 4
    deviation of both eyes to the right side | 4
    unresponsive | 4
    loose stools | 4
    vomiting | 4
    drowsy | 4
    temperature 39.9°C | 4
    oxygen saturation 90% | 4
    blood pressure 72/30 mmHg | 4
    respiratory rate 39/min | 4
    heart rate 220/min | 4
    fluid resuscitation | 4
    high flow oxygen | 4
    loading dose of phenytoin (20 mg/kg) | 4
    electrocardiogram showed sinus tachycardia | 4
    shifted to Intensive Care Unit | 4
    regaining consciousness | 6
    hemodynamically stable | 6
    fully conscious | 9
    normal neurological examination | 9
    shifted out to the pediatric ward | 24
    complete blood count | 24
    serum electrolytes | 24
    blood gases | 24
    serum calcium | 24
    serum magnesium | 24
    glucose levels | 24
    blood culture | 24
    urine culture | 24
    C-reactive protein 0.2 mg/L | 24
    discharged | 72
    phenytoin continued for 3 days after discharge | 72
    phenytoin stopped | 96
    follow-up after 2 months | 1728
    asymptomatic | 1728
    normal neurological examination | 1728
    neuroimaging | 1728
    EEG | 1728

    3 years old | 0
    boy | 0
    admitted | 0
    cough | -48
    cold | -48
    fever | -48
    poor oral intake | -48
    febrile convulsions | -8760
    vomiting | -8760
    cyanosis | -8760
    moderate to high-grade fever | -8760
    deviation of eyes to one side | -8760
    loss of consciousness | -8760
    electroencephalogram (EEG) | -8640
    cerebrospinal fluid studies | -8640
    neuroimaging | -8640
    diagnosis of atypical febrile convulsions | -8640
    no family history of epilepsy | 0
    febrile | 0
    mild congestion in the throat | 0
    symptomatic treatment | 0
    high-grade fever | 4
    vomiting | 4
    bluish discoloration of the extremities | 4
    tachypnea | 4
    deviation of both eyes to the right side | 4
    unresponsive | 4
    loose stools | 4
    vomiting | 4
    drowsy | 4
    temperature 39.9°C | 4
    oxygen saturation 90% | 4
    blood pressure 72/30 mmHg | 4
    respiratory rate 39/min | 4
    heart rate 220/min | 4
    fluid resuscitation | 4
    high flow oxygen | 4
    loading dose of phenytoin (20 mg/kg) | 4
    electrocardiogram showed sinus tachycardia | 4
    shifted to Intensive Care Unit | 4
    regaining consciousness | 6
    hemodynamically stable | 6
    fully conscious | 9
    normal neurological examination | 9
    shifted out to the pediatric ward | 24
    complete blood count | 24
    serum electrolytes | 24
    blood gases | 24
    serum calcium | 24
    serum magnesium | 24
    glucose levels | 24
    blood culture | 24
    urine culture | 24
    C-reactive protein 0.2 mg/L | 24
    discharged | 72
    phenytoin continued for 3 days after discharge | 72
    phenytoin stopped | 96
    follow-up after 2 months | 1728
    asymptomatic | 1728
    normal neurological examination | 1728
    neuroimaging | 1728
    EEG | 1728