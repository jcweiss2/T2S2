30 years old | 0
man | 0
gunshot wounds to the anterior left thoracoabdominal region | -936
gunshot wound to the right back | -936
damage control laparotomy | -936
right nephrectomy | -936
acute kidney injury | -936
haemodialysis | -936
liver injury | -936
bile leak | -936
endoscopic retrograde cholangiogram | -936
common bile duct stent placement | -936
pulmonary embolism | -936
sepsis | -936
prolonged antibiotics | -936
anticoagulation | -936
therapeutic anticoagulation with warfarin | -744
colicky abdominal pain | 0
non-productive cough | 0
Grade III dyspnoea | 0
pyrexia | 0
INR >10 | 0
bilateral pleural effusions | 0
blood products given | 0
empiric broad-spectrum antibiotics | 0
warfarin stopped | 0
respiratory distress | 192
cardiac tamponade | 192
bilateral pleural effusions | 192
cardiomegaly | 192
pericardial effusion | 192
2 cm defect/aneurysm in the lateral right ventricular wall | 192
surgical repair of the right ventricular aneurysm | 216
haemothorax | 192
ejection fraction 45% | 216
bovine pericardial patch | 216
4/0 Prolene suture | 216
focal endarteritis obliterans | 216
therapeutic anticoagulation | 216
follow-up echocardiography | 216
no previous medical history | 0
blood pressure 109/66 mmHg | 0
pulse 95/min | 0
abdomen tender but non-peritonitic | 0
normal chest X-ray | 0
free fluid in the abdomen | 0
arterial blood gas pH 7.18 | 0
lactate 3.5 mmol/L | 0
base excess 5.3 mmol/L | 0
haemoglobin 11 g/dL | 0
HCO3 17 mmol/L | 0
subxiphoid pericardial window | -936
no pericardial effusion | -936
no cardiac injury suspected | -936
normal cardiac examination | -936
normal imaging | -936
first computed tomography unremarkable | -936
intrahepatic collection suggestive of liver abscess | 0
small bilateral pleural effusions | 0
large circumferential pericardial effusion | 192
normal ECG | 192
no ischemic signs | 192
no deep Q waves | 192
Grade 2 pericardial adhesions | 216
cooled to 28°C | 216
bypass perfusion time 132 min | 216
aortic cross-clamp applied | 216
antegrade cold blood cardioplegia | 216
cross-clamp time 41 min | 216
significant bloody pericardial effusion | 216
bile collection in the sub-diaphragmatic area | 216
closed suction drain placed | 216
diaphragmatic defect closed | 216
excised tissue of the RVA 25 x10x3 mm | 216
fibrosis | 216
hemorrhage with organization | 216
haemosiderin deposition | 216
fibrin | 216
dystrophic calcification | 216
granulation tissue | 216
no post-operative complications | 216
satisfactory recovery | 216
no follow-up echocardiography | 216
true aneurysm | 216
false aneurysm | 216
no competing interests | 216
