69 years old | 0  
    man | 0  
    without underlying disease | 0  
    productive cough | -120  
    cold medicine prescribed | -120  
    fever | -24  
    chills | -24  
    breathlessness | -24  
    pain in the right chest wall | -24  
    visited emergency room | 0  
    farmer | 0  
    smoked for 25 years | 0  
    alert | 0  
    blood pressure 90/60 mmHg | 0  
    pulse rate 84/min | 0  
    body temperature 37.1℃ | 0  
    oxygen saturation 79% on room air | 0  
    crackles heard in both lower lung fields | 0  
    arterial blood gas analysis: pH 7.434 | 0  
    arterial blood gas analysis: carbon dioxide partial pressure 34.9 mmHg | 0  
    arterial blood gas analysis: oxygen partial pressure 41.0 mmHg | 0  
    arterial blood gas analysis: bicarbonate 23.6 mmol/L | 0  
    arterial blood gas analysis: oxygen saturation 78.3% | 0  
    white blood cell count 1,710/µL | 0  
    hemoglobin 14.6 g/dL | 0  
    hematocrit 45.1% | 0  
    platelet count 122,000/µL | 0  
    leucopenia | 0  
    no hematologic disease | 0  
    leucopenia recovered spontaneously | 0  
    blood chemistry: urea nitrogen 27 mg/dL | 0  
    blood chemistry: creatinine 1.4 mg/dL |=0  
    blood chemistry: total protein 5.8 g/dL | 0  
    blood chemistry: albumin 3.5 g/dL | 0  
    blood chemistry: aspartate aminotransferase 28 IU/L | 0  
    blood chemistry: alanine aminotransferase 20 IU/L | 0  
    blood chemistry: C-reactive protein 11.40 mg/dL | 0  
    prothrombin time 11.9 seconds | 0  
    activated partial thromboplastin time 34.7 seconds | 0  
    chest X-ray showed haziness in both lower lung fields | 0  
    respiratory distress | 24  
    endotracheal intubation | 24  
    transferred to ICU | 24  
    mechanical ventilator support | 24  
    administered ciprofloxacin | 24  
    administered piperacillin/tazobactam | 24  
    hypoxic despite FiO2 1.0 | 48  
    septic shock despite inotropic agents | 48  
    pneumonia improved progressively | 168  
    suprapubic catheter insertion | 288  
    abdominal pain | 288  
    abdominal computed tomography performed | 288  
    fluid in proximal large intestine | 288  
    reduced contrast enhancement indicating edema in proximal large intestine | 288  
    exploratory laparotomy performed | 288  
    large fluid collection in abdominal cavity | 288  
    necrosis of colon from ileocecal valve to upper rectum | 288  
    no bowel perforation | 288  
    small bowel normal except some inflammatory change | 288  
    subtotal colectomy | 288  
    ileostomy | 288  
    hypoxic damage of bowel during initial hospitalization considered | 288  
    tissue examination during active treatment of septicemia | 288  
    tissue examination during active treatment of acute renal failure | 288  
    colonic infarction due to mucormycosis | 288  
    amphotericin B initiated | 336  
    condition deteriorated | 816  
    died | 816