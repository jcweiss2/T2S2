45 years old | 0
African American male | 0
found unresponsive | -72
supply of K2 within arm's reach | -72
history of depression | -2880
history of anxiety | -2880
history of sleep disorder | -2880
history of hypertension | -2880
history of substance abuse | -2880
elevated blood sugar | -2880
no known history of diabetes | -2880
methadone | -2880
trazodone | -2880
no prior history of neuroleptic agents | -2880
no prior history of serotonin selective reuptake inhibitors | -2880
history of intravenous heroin abuse | -8760
history of inhalational cocaine abuse | -8760
abstinent for the past year | -8760
smoking cannabinoids regularly for 15 years | -131400
using K2 via a bong device twice daily | -504
normal blood pressure (125/81 mmHg) | 0
tachycardia (158 beats/min) | 0
tachypnea (30/min) | 0
high grade temperature (106.5°F) | 0
hypoxia (90% O2 saturation on room air) | 0
obtunded | 0
bilateral pupils equal and reactive to light | 0
normal muscle tone | 0
absence of rigidity | 0
reflexes 1+ and symmetric | 0
no clonus | 0
no focal neurological deficits | 0
regular tachycardia | 0
marked hyperglycemia (Glucose 1,403 mg/dL) | 0
elevated creatinine (3.06 mg/dL) | 0
hypernatremia (Na-160 mmol/L) | 0
hypokalemia (K 2.2 mmol/L) | 0
severe hypophosphatemia (PO4 0.7 mg/dL) | 0
mildly elevated cardiac enzymes (CK 387 U/L, CKMB 1.03 ng/mL, Troponin 0.569 ng/mL) | 0
hepatitis C Ab reactive | 0
HIV Ag/Ab non-reactive | 0
Ab reactivity to hepatitis A and hepatitis B Surface Ag | 0
sinus tachycardia (Heart rate 127/min) | 0
first-degree atrioventricular block | 0
anion gap metabolic acidosis | 0
respiratory acidosis | 0
metabolic alkalosis | 0
hypertriglyceridemia (TG-309 mg/dL) | 0
subarachnoid hemorrhage | 0
possible parenchymal hemorrhage in the left frontal lobe | 0
no soft tissue or bony lesions | 0
focal FLAIR hyper-intense signal | 0
reduction in subarachnoid hemorrhage conspicuity | 24
no evidence of new bleeding | 24
no evidence of trauma | 24
normotensive | 24
normal vasculature on MRA | 24
SC use attributed as cause of intracranial bleeding | 24
no acute neurosurgical intervention | 24
seizure prophylaxis administered | 24
mental status improved | 24
no focal neurological deficit | 24
serial troponin-I levels trended upward | 24
STEMI in leads aVL and I | 24
cardiac risk factors (cigarette smoking, hypertension, diabetes) | 24
denied chest pain | 24
denied shortness of breath | 24
anticoagulation and antiplatelet therapies withheld | 24
hemodynamically stable | 24
mild left ventricular dilation | 24
global hypokinesis | 24
ejection fraction 15% | 24
LV EF improved to 65% | 168
normalization of left ventricle size | 168
no evidence of sepsis | 168
no coronary revascularization | 168
no significant history of alcohol abuse | 168
no apical ballooning on echocardiography | 168
respiratory failure requiring intubation | 168
hyperthermia at admission | 168
no leukocytosis | 168
no bandemia | 168
afebrile for remainder of hospital stay | 168
negative blood cultures | 168
negative sputum cultures | 168
normal urine analysis | 168
normal kidneys on abdominal CT | 168
no source of infection | 168
no cholelithiasis | 168
no cholecystitis | 168
normal chest X-ray on admission | 168
perihilar and bibasilar opacities on day 3 | 72
treated empirically with broad-spectrum antibiotics | 72
changed to ampicillin sulbactam | 72
met SIRS criteria initially | 72
no sources of infection | 72
diagnosed with pneumonia | 72
no SIRS criteria present | 72
normotensive throughout hospitalization | 72
CPK peaked at 301,901 U/L | 336
daily continuous renal replacement therapy | 336
CPK decreased progressively | 336
renal function returned to normal | 336
creatinine 0.95 mg/dL | 336
urine toxicology positive for methadone | 336
negative for cannabinoids | 336
negative for flunitrazepam | 336
negative for gamma hydroxybutarate | 336
recovered entirely to baseline | 504
discharged home | 504
