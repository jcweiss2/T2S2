39 years old | 0
female | 0
ovarian cancer | 0
stage III | 0
TAH with BSO | -432
paclitaxel | -432
carboplatin | -432
melena | -312
hematochezia | -312
abdominal tenderness | -312
rebound tenderness | -312
neutropenia | -312
high fever | -312
tachypnea | -312
hypotension | -312
cyanosis | -312
neutropenic/septic shock | -312
ascending colon perforation | -312
transferred to our hospital | -312
emergent total colectomy | -312
moved to ICU | -312
intubated | -312
alert | -312
oriented | -312
difficulty in weaning from mechanical ventilation | -312
severe tachypnea | -312
labored breathing | -312
sedated with midazolam | -288
neutropenia did not improve | -288
ANC less than 50/µl | -288
chemotherapy induced neutropenia | -288
sepsis suspected | -288
G-CSF administered | -288
antibiotics administered | -288
midazolam stopped | -240
extubated | -240
dyspnea | -240
deteriorating levels of consciousness | -240
reintubation | -240
brain CT | -240
EEG performed | -240
no abnormal findings on brain CT | -240
no abnormal findings on EEG | -240
neurologic status did not improve | -216
partial seizure | -216
generalized tonic-clonic seizure | -216
seizure controlled with midazolam | -216
seizure controlled with ativan | -216
seizure controlled with phenytoin | -216
diffuse brain swelling | -216
severe diffuse cerebral dysfunction on EEG | -216
severe hyperammonemia | -216
arterial blood gas analysis showed respiratory alkalosis | -216
arterial blood gas analysis showed metabolic alkalosis | -216
electrolytes unremarkable | -216
liver panel unremarkable | -216
CRRT administered | -216
follow-up ammonia level 1,356 µg/dl | -216
sodium benzoate administered | -216
mannitol administered | -216
recurrent episodes of GTC seizure | -216
status epilepticus | -216
midazolam administered | -216
phenytoin administered | -216
further partial seizures | -216
desaturation | -216
hypotension | -216
died | -168
