25 years old|0
woman|0
low back pain|0
intravenous drug use|0
hypotension|0
hypoxemic respiratory failure|0
intubation|0
transthoracic echocardiography|0
large mobile tricuspid vegetations|0
severe tricuspid regurgitation|0
chest radiograph|0
extensive bilateral patchy opacifications|0
recurrent episodes of pulseless electrical activity|0
veno7arterial extracorporeal membrane oxygenation cannulation|0
right femoral vein|0
right femoral artery|0
antegrade catheter|0
distal limb perfusion|0
refractory hypoxemia|0
temperature 97.5 °F|0
heart rate 74 beats/min|0
sinus rhythm|0
blood pressure 88/56 mm Hg|0
norepinephrine 5 μg/min|0
oxygen saturation 84%|0
6 L/min VA7ECMO|0
maximal oxygenation on ventilator|0
right radial arterial blood gas analysis|0
PaO2 of 44 mm Hg|0
blood cultures grew methicillin-sensitive Staphylococcus aureus|0
transesophageal echocardiography|0
mildly reduced biventricular systolic function|0
multiple tricuspid valve vegetations|0
valve perforation|0
severe TR|0
no other vegetations|0
no intracardiac shunt|0
computed tomography|0
extensive lung consolidative and cavitary opacities|0
small pleural effusions|0
sacroiliitis|0
no intracranial process|0
percutaneous aspiration strategy|0
severe right-side endocarditis|0
differential hypoxemia|0
preserved cardiac output|0
poorly oxygenated blood|0
north-south syndrome|0
Harlequin syndrome|0
maximization of ECMO flows|0
pulmonary optimization|0
ventilator adjustments|0
airway clearance maneuvers|0
targeted therapy|0
severe ongoing airway bleeding|0
purulent mucous|0
substantial septic pulmonary emboli|0
transition to veno7arterial7venous ECMO|0
introduction of additional return cannula|0
Y-configuration|0
improved peripheral oxygenation|0
hemodynamic compromise|0
venous access|0
serial dilations|0
ECMO flows reduced|0
de-airing techniques|0
occluder device|0
Hoffman clamp|0
inotropic support|0
cardiac output|0
VA7ECMO weaning method|0
multidisciplinary meeting|0
heart team meeting|0
cardiology|0
cardiothoracic surgery|0
cardiac anesthesia|0
pulmonary|0
nursing|0
medical ethics|0
not a surgical candidate|0
severe lung injury|0
percutaneous aspiration of tricuspid vegetations|0
trivial echodensity|0
stable severe TR|0
veno-venous extracorporeal circuit|0
filter and pump|0
reinfusion of blood|0
left internal jugular|0
left femoral vein|0
therapeutic anticoagulation|0
clamping of arterial limb|0
hemodynamics on VV bypass|0
low-dose vasopressor support|0
cannulation strategies for VV7ECMO|0
drainage cannula|0
return cannula|0
femoral vein|0
right internal jugular vein|0
IVC7RA junction|0
SVC7RA junction|0
femoral-femoral VV7ECMO|0
single dual-lumen ECMO cannula|0
ProtekDuo|0
dual-lumen cannula|0
main pulmonary artery|0
right ventricle decompression|0
hemodynamically stable|0
impaired respiratory gas exchange|0
transition to VV7ECMO|0
dual lumen catheter|0
ongoing hypoxemia|0
recirculation|0
membrane dysfunction|0
cannula malposition|0
membrane lung shunting|0
increased sedation|0
calcium channel blockers|0
beta-blockers|0
negative inotropic agents|0
right ventricular dysfunction|0
second venous drainage cannula|0
second parallel VV7ECMO circuit|0
esmolol infusion|0
high cardiac output|0
prolonged course of intravenous antibiotics|0
MSSA infection|0
bronchopleural fistula|0
empyema necessitans|0
video-assisted thorascopic surgery|0
Eloesser flap|0
improved airway bleeding|0
improved pleural disease|0
decannulation from VV7ECMO|0
preserved left ventricular function|0
dilated right ventricle|0
normal systolic function|0
persistent severe TR|0
small vegetation|0
prolonged critical illness|0
discharged|0
intensive physical therapy|0
ongoing care|0
no dyspnea|0
no heart failure symptoms|0
