37 years old | 0
female | 0
admitted to the hospital | 0
parity 3 | 0
gestation 2 | 0
vaginal delivery | -96
lateral episiotomy | -96
spontaneous vaginal delivery of twins | -96
serologic testing of HIV | -96
serologic testing of hepatitis | -96
vaginal swabs | -96
urine culture | -96
discharged after 24 h | -72
nonspecific abdominal pain | 0
septic shock | 0
axillary temperature 36 °C | 0
blood pressure 80/30 mmHg | 0
tachycardia 130/min | 0
marbling | 0
cold limbs | 0
abdominal ultrasound | 0
free intra-abdominal fluid | 0
fluid resuscitation | 0
catecholamine | 0
noradrenaline | 0
tachypneic | 0
respiratory rate 30 cycle/min | 0
unspecific bowel infection | 0
broad-spectrum antimicrobial treatment | 0
imipenem | 0
amikacin | 0
teicoplanin | 0
hemoglobin level 9.2 g/dL | 0
leukocytes 1540 × 10 [3]/μL | 0
platelet count 104000/μL | 0
C-reactive protein 340 mg/dL | 0
creatinine 1.92 mg/dL | 0
albumin 1.2 g/dL | 0
cytolysis | 0
ALT 120 UI/L | 0
AST 146 UI/L | 0
cholestasis | 0
blood gas | 0
metabolic acidosis | 0
pH 7.12 | 0
arterial lactate levels 8.9 mmol/L | 0
SOFA score 9 | 0
emergency exploratory laparotomy | 2
purulent fluid | 2
global venous congestion | 2
inspection of the bladder | 2
inspection of the uterus | 2
inspection of the adnexa | 2
inspection of the bowel | 2
lavage of the peritoneal cavity | 2
pelvic drain | 2
heparin | 2
CT scan of the abdomen | 4
intraperitoneal free fluid | 4
paralytic ileus | 4
no sign of arterial or venous thrombosis | 4
fluid culture | 6
blood culture | 6
group A streptococci | 6
septic shock | 6
multiorgan failure | 6
disseminated intravascular coagulation | 6
death | 12