43 years old | 0
man | 0
pedestrian accident | 0
admitted to the hospital | 0
comatose | 0
Glasgow coma score of 3 | 0
nonreactive pupils 5 mm in diameter | 0
ventilated | 0
hemodynamically stable condition | 0
bilateral otorrhea | 0
rhinorrhea | 0
bruising in face | 0
bruising in jaw | 0
bruising in right side of the scalp | 0
diffuse brain injury | 0
severe cerebral swelling | 0
right-side acute subdural hemorrhage | 0
ring fracture around the foramen magnum | 0
clivus fracture | 0
petrous temporal bones fracture | 0
posterior part of the foramen magnum fracture | 0
no atlanto1-occipital dislocation | 0
cervical spine intact | 0
admitted to the neurosurgical intensive care unit | 0
no subsequent neurological changes | 0
brain death suspected | 0
healthy before the accident | -672
coma | 0
Glasgow coma scale score of 3 | 0
fixed, nonreactive pupils 6 mm in diameter | 0
no signs of brain stem activity | 0
vital signs stable | 0
swelling of the brain stem | 648
swelling of the cerebellum | 648
transtentorial herniation | 648
foraminal herniation | 648
pontomedullary laceration | 648
fully comatose | 0
pneumonia | 816
sepsis | 816
died | 816
ring fracture | 0
sudden heart arrest | 0
cerebrospinal fluid rhinorrhea | 0
cerebrospinal fluid otorrhea | 0
no combined injury | 0
severe cerebral swelling |5 0
no atlanto-occipital dislocation | 0
