Here is the table of events and timestamps:

70 years old | 0
male | 0
emergency esophageal diversion | 0
injury to the cervical esophagus | 0
esophageal diversion | 0
retrosternal GPU procedure | -168
postoperative anastomotic leakage | -168
endoscopy | -168
fully covered esophageal stent | -168
discharged | -168
local cervical infection | -84
sepsis | -84
transferred to the intensive care unit | -84
antibiotic treatment | -84
endoscopy | -84
dislocated stent | -84
pus evacuation and debridement | -84
fully covered self-expanding metal stent | -84
percutaneous jejunal feeding catheter | -84
re-endoscopy | -84
slippage of the stent | -84
EVT | -84
EsoSponge system | -84
jugular and cervical phlegmon resolved | -56
repeated endoscopic balloon dilatation | -56
subtotal esophageal resection and reconstruction | 0
free-jejunal graft interposition | 0
partial sternotomy | 0
laparotomy | 0
jejunal segment harvested | 0
cervical anastomosis | 0
upper mediastinal gastro-jejunostomy | 0
abdominal reconstruction | 0
oral alimentation | 24
speech therapy | 24
anastomotic healing | 24
transferred to a rehabilitation clinic | 24