61 years old | 0
male | 0
non-Hodgkin’s lymphoma | -10080
prior radiation therapy | -10080
coronary artery disease | -10080
coronary artery bypass graft | -10080
mechanical aortic valve replacement | -10080
severe bicuspid aortic valve stenosis | -10080
admitted to the hospital | 0
fever | -72
malaise | -72
respiratory distress | -72
broad-spectrum intravenous antibiotics | -72
sepsis | -72
intubated | -72
respiratory failure | -72
methicillin-sensitive Staphylococcus aureus | -72
transesophageal echocardiogram | -72
vegetation on the mechanical aortic valve | -72
prosthetic endocarditis | -72
intravenous oxacillin | -72
gentamicin | -72
rifampin | -72
pulseless electrical activity cardiac arrest | -144
complete heart block | -144
external MRI-compatible pacemaker | -144
right ventricle MRI-compatible active-fixation lead | -144
left subclavian approach | -144
stenosis of the internal jugular veins | -144
computed tomography of the head | -138
multifocal bilateral infarcts | -138
small areas of adjacent parenchymal and subarachnoid hemorrhage | -138
persistent ventilator requirement | -120
left pneumothorax | -120
chest tube placement | -120
progressive renal injury | -120
acute tubular necrosis | -120
transferred to our institution | -120
intubated | -120
sedated | -120
corneal and gag reflexes were present | -120
grimaced in response to upper extremity noxious stimuli | -120
no response to lower extremity noxious stimuli | -120
white blood count of 22,700/μL | -120
hemoglobin 9.4 g/dL | -120
platelets 402,000/μL | -120
creatinine 3.2 mg/dL | -120
limited transthoracic echocardiogram | -120
aortic valve vegetation | -120
trace aortic regurgitation | -120
brain MRI | -108
septic emboli | -108
developing brain abscess | -108
contrast CT imaging | -108
renal insufficiency | -108
noncontrast CT | -108
Magnetic Resonance Safety Officer | -108
MR Medical Director | -108
1.5 T MR scanner | -108
transmit-receive head coil | -108
normal mode | -108
repositioning of the generator | -108
insulating the generator | -108
gauze pads | -108
transparent film dressing | -108
complete heart block | -108
ventricular escape | -108
pre-MRI impedance | -108
threshold values | -108
pacemaker MRI mode | -108
VOO at 80 beats per minute | -108
pacing output of 5.0 V at 1.0 ms | -108
transcutaneous pacing pads | -108
external defibrillator | -108
intensive care nurse | -108
continuous telemetry | -108
pulse oximetry | -108
35 minutes of scanning | -108
post-MRI impedance | -72
thresholds | -72
battery capacity | -72
chest roentgenograph | -72
lead migration | -72
brain MRI images | -72
bilateral multifocal infarcts | -72
septic emboli | -72
brain abscess | -72
cardiac CT | -48
aortic root abscess | -48
benzodiazepine | -48
neuromuscular blockade | -48
breath-holding | -48
VOO at 70 beats per minute | -48
motion artifact | -48
large hypoattenuated mass | -48
vegetation | -48
thickening of the mitral-aortic intervalvular fibrosa | -48
perivalvular involvement | -48
no abscess | -48
lead position | -48
right ventricular apex | -48
cardiac surgery | -24
operative mortality risk | -24
surgical intervention | -24
palliative care | -24
comfort-oriented care | -24
died | 0