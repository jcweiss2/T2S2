56 years old| 0
male | 0
breathlessness on exertion | -17520
breathlessness at rest | -17520
prolonged cough | -17520
bloody sputum production | -17520
hoarseness | -17520
decline in performance impact | -17520
reduced tolerance to physical activity | -17520
breathlessness | -17520
chronic bronchitis | -17520
antibacterial therapy | -17520
mucolytic therapy | -17520
local therapy | -17520
admitted | 0
significant decrease of blood oxygenation | 0
NYHA III-IV condition | 0
stridor | 0
respiratory distress | 0
preoperative chest CT | -24
giant ascending aorta | -24
aortic arch | -24
thoracic aorta partially-thrombosed ampullary false aneurysm | -24
left main bronchus compression | -24
left pulmonary artery compression | -24
trachea compression | -24
left pulmonary veins compression | -24
esophagus compression | -24
azygos vein compression | -24
recurrent pneumonia | -24
trachea drainage tube disorder | -24
multivessel coronary artery disease | -24
surgery performed as emergency | 0
cardiopulmonary bypass | 0
right subclavian artery cannulation | 0
central venous cannulation | 0
supra-bifurcation compression of the trachea | 0
compression of the left main bronchus | 0
tracheal intubation using bronchoscopy | 0
complete compression of the left main bronchus | 0
right lung ventilation | 0
distal anastomoses of the coronary artery bypass grafting | 0
target temperature 26°C | 0
ascending aorta mobilised | 0
aneurysmal sac separated from pulmonary artery branches | 0
ascending aorta transected | 0
blood antegrade cardioplegia | 0
brachiocephalic trunk clamped | 0
visceral arrest | 0
monohemispheral perfusion of the brain | 0
aneurysmal sac opened | 0
intimal rupture | 0
massive thrombotic masses | 0
sac excised | 0
aneurysm bed sanitized | 0
affected aorta cut off | 0
aorta-tracheal fistula found | 0
temporarily damped with antiseptic napkin | 0
total replacement of the aortic arch | 0
synthetic multi-branch prosthesis | 0
supracoronary replacement of ascending aorta | 0
proximal anastomosis with prosthesis | 0
coronary arteries bypass grafts | 0
trachea exposed | 0
suture repair of the postero-lateral wall defect | 0
tightness control using bronchoscopy | 0
decompression of the airways | 0
endotracheal tube repositioned | 0
left lung included | 0
extubated | 48
observation in intensive care unit | 48
bronchoscopy control for tightness | 48
bronchoscopy control for patency | 48
discharged | 336
satisfactory echocardiography | 336
satisfactory laboratory tests | 336
no data for respiratory failure | 336
no data for heart failure | 336
no data for coronary failure | 336
dynamic CT | 336
no infiltrative changes in the lungs | 336
no infiltrative changes in the mediastinum | 336
histological examination | 336
atherosclerosis | 336
thinning of aortic wall tissue | 336
inflammation of aortic wall tissue | 336
NYHA I | 8760
CT follow-up | 8760
no special features in aortic arch reconstruction area | 8760
patency of the trachea restored | 8760
patency of the main bronchus restored | 8760
