66 years old | 0
    female | 0
    presented with diffuse pruritus | -432
    presented with erythroderma | -432
    biopsy revealed atypical cells | -432
    flow cytometry showed abnormal CD3+ CD4+ CD7− CD26− T-cell clone | -432
    hematopathology showed Sézary cell count of 2312 | -432
    positron emission tomography scan showed bilateral lymphadenopathy | -432
    stage IVA1 (T4NxM0B2) Sézary syndrome | -432
    uncontrolled hypertension | 0
    type 2 diabetes | 0
    end-stage renal disease | 0
    prescribed extracorporeal photopheresis | -432
    prescribed bexarotene | -432
    lost to follow-up | -432
    pruritus worsened | -432
    Sézary count climbed to 11,132 | -432
    April 2020 SARS-CoV-2 infection | -24
    shortness of breath | -24
    afebrile | -24
    recovered fully without medication | -24
    Sézary count dropped to 6494 | 168
    July 2020 admission | 0
    severe COVID-19 | 0
    shortness of breath | 0
    chills | 0
    fever (38.5 °C) | 0
    hypoxemia (70% O2 saturation) | 0
    protracted 25-day stay | 0
    multiple ICU admissions | 0
    received dexamethasone | 0
    received empiric antibiotics | 0
    false-positive blood culture | 0
    lymphocyte count began to decrease on hospital day 14 | 336
    discharge with absolute lymphocyte count of 1900 | 600
    September 2020 clinic return | 2160
    Sézary count dropped to 936 | 2160
    began romidepsin therapy | 2160
    October 2020 improved pruritus | 2880
    resolved erythroderma | 2880
    resolved lymphadenopathy | 2880
    Sézary counts dropped to 389 | 2880
    November admission | 3384
    severe COVID-19 | 3384
    developed encephalopathy | 3384
    hypotension | 3384
    cardiac arrest | 3384
    death | 3384
    papulonodular rash | -432
    lymphadenopathy | -432
    diffuse pruritus | -432
    erythroderma | -432
    CD4:CD8 ratio 6 | -432
    CD4:CD8 ratio 22.5 | -432
    CD4:CD8 ratio 23 | 168
    CD4:CD8 ratio 6.3 | 2880
    improved pruritus | 2880
    continued papulonodular rash | 2880
    resolved lymphadenopathy | 2880
    resolved erythroderma | 2880
    no SS treatment until September 2020 | 2160
    denied SS treatment during July 2020 admission | 0
    denied chest pain | 0
    no shortness of breath in April 2020 | -24
    negative COVID-19 test in July readmission | 0
    no fever in April 2020 | -24
    negative blood culture during July admission | 0