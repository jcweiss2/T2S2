27 years old | 0
male | 0
admitted to the psychiatric department | 0
acute psychiatric syndrome | 0
personality and behavioral change | 0
friendly | 0
focused attention | 0
clear consciousness | 0
responded slowly to questions | 0
emotional instability | 0
interruption of thinking | 0
thinking burst | 0
absence of hallucination | 0
absence of delusion | 0
absence of impulsive aggression | 0
psychotropic drugs | 0
rigidity | 7
transferred to neurology department | 12
suspected viral encephalitis | 12
neurological impairment | 12
abnormal movements | 12
tachycardia | 12
status epilepticus | 12
insomnia | 12
confusion of consciousness | 12
memory deficits | 12
absence of fever | 12
electroencephalogram (EEG) | 12
diffuse or general slowing | 12
magnetic resonance imaging (MRI) of the brain | 12
no abnormal changes | 12
cerebrospinal fluid (CSF) analysis | 12
mild elevations of the protein level | 12
elevations of the karyocyte count | 12
normal glucose level | 12
antibody against NR1 heteromeric NMDAR detected | 12
comprehensive tumor screening | 12
no tumors or inflammatory lesions detected | 12
diagnosed with ANMDARE | 12
treated with anti-epileptic drugs | 12
corticosteroids | 12
intravenous immunoglobulin (IVIG) | 12
improved and discharged | 24
new hyperpyrexia | -24
dyspnea | -24
severe status epilepticus | -24
decreased level of consciousness | -24
convulsion of the limbs | -24
admitted to the emergency intensive care unit (EICU) | -24
supplemental oxygen | -24
perspiration | -24
cutaneous pallor | -24
mild tachypnea | -24
severe hypoxemia | -24
good air entrance bilaterally | -24
scattered to diffuse crackles and rhonchi | -24
elevated serum C-reactive protein | -24
elevated procalcitonin (PCT) | -24
acute lung inflammation on CT | -24
abnormal CSF | -24
positive anti-NMDAR antibodies | -24
negative Herpes simplex virus (HSV) DNA PCR | -24
Acinetobacter baumanii in sputum culture | -24
relapse of anti-NMDAR encephalitis | -24
pneumonia caused by acinetobacter baumannii | -24
treated with steroid and IVIG pulse therapy | -24
antibacterial agents | -24
supportive therapies | -24
gradually recovered | 0
mild psychiatric sequelae | 0