52 years old | 0
female | 0
admitted to the hospital | 0
fever | -240
cough | -240
breathlessness | -240
progressive dyspnea | -240
respiratory distress | -240
decrease urine output | -240
no abdominal pain | -240
no dysuria | -240
no trauma | -240
no recent use of non-steroidal anti-inflammatory medication | -240
breathless | 0
blood pressure 150/90 mmHg | 0
temperature 40°C | 0
respiratory rate of 30 breaths/min | 0
heart rate of 100 bpm | 0
hemoglobin 10.3 g/l | 0
total white cell count 9.88 × 10^3/μl | 0
differential count: 74% neutrophils, 20% lymphocytes, 4% monocytes and 2% eosinophils | 0
platelet count 211 × 10^3/μl | 0
serum creatinine 10.8 mg/dl | 0
sodium 138 mEq/l | 0
potassium 5.3 mEq/l | 0
blood urea 76 mg/dl | 0
blood glucose 72 mg/dl | 0
normal sized kidneys with hyper reflective cortex | 0
negative serological tests for malaria, leptospirosis, dengue and viral hepatitis | 0
sterile blood, urine and sputum cultures | 0
proteinuria | 0
hematuria | 0
two to five fine granular casts | 0
oseltamivir treatment | 0
antibiotic treatment | 0
fluid replacement | 0
dialysis | 0
peritoneal dialysis | 0
intermittent hemodialysis | 0
renal biopsy | 24
mesangial proliferative glomerulonephritis | 24
acute tubule interstitial nephritis | 24
methyl prednisolone treatment | 48
oral prednisolone treatment | 48
discharged | 168
SCr 1.5 mg/dl | 168
SCr 1 mg/dl at 1 month follow-up | 720