48 years old | 0
man | 0
admitted to the Proctology Department | 0
medical history of syphilis | 0
no treatment due to penicillin anaphylaxis | 0
TRUST value 1:1 | 0
treated with etimicin | -48
treated with ornidazole | -48
incision and drainage for perianal abscess | 0
neck pain | 1
dizziness | 1
chest pressure | 1
high blood pressure 160/90 mmHg | 1
fever 40°C | 2
decreased blood pressure 80/50 mmHg | 2
neutrophilic leukocytosis | 2
procalcitonin level 66.9 ng/mL | 2
temperature dropped to 36.8°C | 2
transferred to ICU | 2
treated with intravenous imipenem-cilastatin | 48
treated with dopamine | 48
worsening neutrophilic leukocytosis | 72
procalcitonin > 200 ng/mL | 72
developed MODS | 96
abscess culture revealed Neisseria gonorrhoeae | 96
abscess culture revealed Staphylococcus haemolyticus | 96
blood cultures revealed R. mannitolilytica | 96
changed to ceftriaxone | 96
changed to levofloxacin | 96
repeat blood cultures no bacterial growth | 192
incision wound healed | 192
satisfactory recovery | 192
6-month follow-up | 4320
no complications | 4320
