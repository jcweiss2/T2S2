history of arterial hypertension | -1000
history of obesity | -1000
fever | -336
mild cough | -336
rhinitis | -336
admission | 0
hypotension | 0
asthenia | 0
alert | 0
oriented | 0
cooperative | 0
asthenic | 0
blood pressure 85/55 mmHg | 0
heart rate 120 bpm | 0
arterial oxygen saturation 85% | 0
fever with body temperature 38.3 C° | 0
femoral central venous catheter positioned | 0
sinus tachycardia | 0
diffuse low voltages | 0
absence of significant repolarization abnormalities | 0
neutrophilic leukocytosis | 0
C-reactive protein elevation | 0
Procalcitonin elevation | 0
elevated high sensitivity Troponin | 0
elevated brain natriuretic peptide | 0
elevated creatinine | 0
elevated transaminases | 0
elevated total bilirubin | 0
negative RT-PCR nasopharyngeal swab for COVID-19 | 0
high COVID-19 IgM antibody | 0
normal left ventricular cavitary dimensions | 0
diffuse LV parietal thickening | 0
severely reduced LV global systolic function | 0
grade II LV diastolic dysfunction | 0
normal cavitary dimensions | 0
reduced global right ventricular systolic function | 0
dilated inferior vena cava | 0
right ventricular systolic pressure 41 mmHg | 0
absence of hemodynamically significant valvulopathy | 0
slight pericardial effusion | 0
broad-spectrum antibiotic therapy started | 0
crystalloid hydration started | 0
nasal cannula ventilatory therapy started | 0
norepinephrine therapy started | 0
poor hemodynamic response to norepinephrine | 12
levosimendan therapy started | 12
blood pressure increased to 100/60 mmHg | 12
heart rate decreased to 110 bpm | 12
further hemodynamic improvement | 24
blood pressure 125/70 mmHg | 24
heart rate 95 bpm | 24
diuresis 1800 ml | 24
improvement of systolic performance indices | 24
improvement of LV diastolic function | 24
removal of central venous catheter | 48
negative culture of CVC tip | 48
cardiac magnetic resonance imaging performed | 72
endomyocardial biopsy performed | 96
discharge | 504
normal laboratory findings at discharge | 504
normal electrocardiographic findings at discharge | 504
normal echocardiographic findings at discharge | 504
normal TTE at 1 month after discharge | 744
normal TTE at 3 months after discharge | 1104