93 years old | 0
male | 0
admitted to the hospital | 0
syncopal episode | 0
coronary heart disease | -6720
percutaneous coronary intervention | -144
stent implantation | -144
dual antiplatelet therapy | -144
atrioventricular pacemaker implantation | -10080
ventricular pacemaker lead replacement | 0
LBB pacing lead implantation | 0
severe fall in blood pressure | 1
pallor | 1
signs of hypoperfusion | 1
shock | 1
inverted T waves | 1
reduced left ventricular function | 1
apical dyskinesis | 1
LV outflow tract obstruction | 1
moderate-to-severe mitral regurgitation | 1
cardiac catheterization | 2
no obstruction in coronary arteries | 2
apical ballooning | 2
basal hyperkinesia | 2
intra-aortic balloon pump | 2
intensive care unit | 2
inotropes avoided | 2
dobutamine avoided | 2
improved hemodynamics | 120
IABP removed | 120
complete resolution of LVOT obstruction | 120
apical ballooning resolved | 120
LV function recovered | 120
EF of 50% | 504
regression of inverted T waves | 504
septic shock | 840
ventilation-associated pneumonia | 840
death | 840
ventricular noise reversion | -1
asystole periods | -1
pacemaker inhibition | -1
ventricular oversensing | -1
Holter monitoring | -1
arterial hypertension | 0
right bundle branch block | 0 
right ventricular lead extraction | 0 
new LBB pacing lead placement | 0 
cardiogenic shock management | 1 
cardiac marker levels normal | 0 
echocardiography normal | 0 
ejection fraction 63% | 0 
electrocardiogram normal | 0 
chest radiography normal | 0 
blood pressure 112/68 mm Hg | 0 
heart rate 60 beats/min | 0 
physical examination normal | 0 
atrial and ventricular stimulation | 0 
DDD mode | 0 
heart rate 60 beats/min | 0 
inotropes started | 48 
LVOT obstruction reduced | 48 
basal hyperkinesia reduced | 48 
apical ballooning reduced | 48 
EF improved | 120 
inotropes effective | 120 
IABP support | 2 
ICU support | 2 
septic shock treatment | 840 
ventilation-associated pneumonia treatment | 840 
cardiac function partially recovered | 504 
pacing parameters stable | 504 
capture threshold stable | 504 
sensing stable | 504 
R wave stable | 504 
ventricular function improved | 504 
inotropes effective | 504 
EF 50% | 504 
inverted T waves regressed | 504 
LBB pacing effective | 504 
physiological ventricular activation | 504 
dyssynchrony reduced | 504 
LV dysfunction improved | 504 
resynchronization therapy effective | 504 
perioperative care crucial | 0 
prompt recognition crucial | 0 
management crucial | 0 
Takotsubo cardiomyopathy diagnosed | 1 
TCM triggered by LBB pacing | 1 
TCM rare in older men | 1 
TCM severe course | 1 
heart failure | 1 
cardiogenic shock | 1 
intensive care unit support | 2 
left ventricular outflow tract obstruction | 1 
inotropes avoided | 2 
basal hyperkinesia | 1 
apical ballooning | 1 
inotropes contraindicated | 2 
inotropes worsen obstruction | 2 
IVPG increased | 2 
hemodynamic parameters deteriorated | 2 
clinical teams aware | 0 
surgical teams aware | 0 
prompt therapeutic management | 2 
unique clinical characteristics | 2 
unique hemodynamic characteristics | 2 
LBB pacing modality | 0 
His bundle pacing modality | 0 
physiological ventricular activation | 0 
clinical indications growing | 0 
complications relatively unknown | 0 
LBB pacing elicits TCM | 1 
perioperative care crucial | 0 
prompt recognition crucial | 0 
management crucial | 0 
TCM incidence increased | 0 
conventional RV pacing triggers TCM | 0 
LBB pacing triggers TCM | 0 
older men rare | 0 
severe course | 0 
heart failure | 0 
cardiogenic shock | 0 
intensive care unit support | 0 
left ventricular outflow tract obstruction | 0 
inotropes avoided | 0 
basal hyperkinesia | 0 
apical ballooning | 0 
inotropes contraindicated | 0 
inotropes worsen obstruction | 0 
IVPG increased | 0 
hemodynamic parameters deteriorated | 0 
clinical teams aware | 0 
surgical teams aware | 0 
prompt therapeutic management | 0 
unique clinical characteristics | 0 
unique hemodynamic characteristics | 0 
LBB pacing modality | 0 
His bundle pacing modality | 0 
physiological ventricular activation | 0 
clinical indications growing | 0 
complications relatively unknown | 0 
LBB pacing elicits TCM | 0 
perioperative care crucial | 0 
prompt recognition crucial | 0 
management crucial | 0