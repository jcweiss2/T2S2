72 years old | 0
woman | 0
admitted for fever | 0
pain in bilateral big toes | 0
no history of trauma | 0
no insect bites recently | 0
episodes happen twice a year | 0
resolves spontaneously | 0
Traditional Chinese Medicine use | 0
negative drug toxicology screen | 0
no diagnosis of gout | 0
no autoimmune problem | 0
negative vasculitis screen | 0
borderline positive anti-nuclear antibody | 0
no risk factors for peripheral vascular disease | 0
pain on bilateral big toes | 0
bilateral podagra | 0
minimal swelling | 0
full range of motion | 0
pulses well felt | 0
admitted to Medical Intensive Care Unit | 0
streptococcal septicaemia | 0
Streptococcus pneumoniae in blood culture | 0
broad spectrum antibiotics started | 0
hypotension 60/40 mmHg | 0
urine output <20 ml/h | 0
no response to fluid replacement | 0
dopamine use up to 18 mcg/kg/min | 0
noradrenaline use up to 0.5 mcg/kg/min | 24
vital signs normalized | 0
dusky extremities | 0
marked livedo reticularis | 48
ecchymosis | 120
mottled skin | 120
necrotic terminal digits | 120
necrotic tip of nose | 120
dry gangrene signs | 120
ecchymotic bullae over bilateral lower limbs | 168
plantar gangrene | 168
non-palpable dorsalis pedis pulses | 168
non-palpable posterior tibial pulses | 168
ecchymotic bullae over bilateral hands | 168
ecchymotic bullae over forearms | 168
non-palpable radial pulses | 168
dry gangrene involved all digits | 168
microvascular spasm diagnosis | 168
no pulsations in gangrenous extremities | 168
arterial occlusion test revealed moderate calcification | 168
referral to plastic surgery | 168
dry gangrene demarcation plan | 168
dry gangrene progressed to bilateral ankles | 720
dry gangrene progressed to wrists | 720
demarcation up to upper forearms | 720
demarcation up to mid-shin left lower limb | 720
demarcation up to upper shin right lower limb | 720
elective re-admission two months later | 1440
four limb amputations | 1440
bilateral below knee amputations | 1440
bilateral above elbow amputations | 1440
smooth recovery post-operatively | 1440
rehabilitation started | 1440
ambulatory with prosthesis | 52560
lower limb prosthesis installed | 4320
upper limb prosthesis utilization | 52560
