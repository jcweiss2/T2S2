70 years old | 0
male | 0
farmer | 0
admitted to the hospital | 0
high-grade fever | -120
generalized body ache | -120
headache | -120
altered sensorium | -24
joint pains | -120
epigastric pain | -120
no comorbidities | 0
no drug addiction | 0
no intoxication | 0
inguinal lymphadenopathy | 0
mild generalized rash | 0
no eschar | 0
hemodynamically stable | 0
disoriented | 0
no focal neurological deficit | 0
no neck rigidity | 0
acute febrile illness | 0
undifferentiated fever | 0
workup for tropical infections | 0
malaria test negative | 0
dengue test negative | 0
typhoid test negative | 0
leptospira test negative | 0
scrub typhus antigen card positive | 0
scrub immunoglobulin M positive | 0
diagnosis of scrub typhus | 0
blood cultures sterile | 0
body fluid cultures sterile | 0
leukocytosis | 0
mild hyperbilirubinemia | 0
transaminitis | 0
slightly raised international normalized ratio | 0
hepatitis B antigen negative | 0
hepatitis C antibody negative | 0
mild fatty infiltration of the liver | 0
tablet doxycycline 100 mg twice daily | 0
defervescence | 48
improved orientation | 48
weakness of both lower limbs | 96
weakness progressed to upper limbs | 96
deep tendon reflexes absent | 96
plantar responses flexor | 96
bladder incontinence | 96
no bowel incontinence | 96
breathing difficulty | 96
respiratory distress | 96
single breath count 10 | 96
respiratory acidosis | 96
intubated | 96
mechanical ventilation | 96
MRI of the brain normal | 96
MRI of the cervical spine normal | 96
nerve conduction velocity showed motor sensory demyelinating polyneuropathy | 96
diagnosis of GBS | 96
cerebrospinal fluid analysis | 96
albuminocytologic dissociation not present | 96
intravenous immunoglobulin therapy | 96
tablet rifampicin 600 mg twice daily | 96
improvement in weakness | 144
improvement in respiratory parameters | 144
weaned off ventilator | 240
extubated | 240
oral feeding started | 240
aggressive limb and chest physiotherapy | 240
shifted out of ICU | 240
discharged from hospital | 672
full neurological recovery | 672