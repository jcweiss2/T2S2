Here is the table of events and timestamps:

54 years old | 0
male | 0
pre-syncope | -4
syncope | -4
left-sided chest tightness | -4
generalized fatigue | -4
weight loss | -4
admitted to the hospital | 0
weight | 0
blood pressure | 0
cardiac examination | 0
respiratory examination | 0
diffuse erythematous rash | 0
electrocardiography | 0
normal sinus rhythm | 0
raised troponin concentration | 0
eosinophil count | 0
referred to cardiology | 0
myocarditis | 0
cardiac magnetic resonance imaging | 0
eosinophilic myocarditis | 0
coronary angiography | 0
no evidence of coronary artery disease | 0
skin biopsy | 0
eczematous changes | 0
bone marrow biopsy | 0
no increase in eosinophils | 0
axillary lymph node biopsy | 0
T-cell lymphoma | 0
improved clinically | 0
discharged | 0
prescribed edoxaban | 0
prescribed prednisolone | 0
follow-up in the rheumatology clinic | 0
missed follow-up | 72
neck swelling | 72
urgent admission to hospital | 72
rise in eosinophil count | 72
increased dose of prednisolone | 72
computed tomography of the neck | 72
lymphadenopathy | 72
T-cell lymphoma confirmed | 72
course of chemotherapy with cyclophosphamide | 72
sepsis secondary to cholecystitis | 72
new onset of seizures | 72
reduction in consciousness | 72
Glasgow Coma Scale 9/15 | 72
head CT | 72
multiple bilateral acute infarctions | 72
investigations to identify the source of the infarcts | 72
history of hepatitis B | -4
history of asthma | -4
history of intravenous drug use | -4
history of excessive alcohol use | -4
apical tear | 72
intramural myocardial tear | 72
small apical cavity | 72
mobile structures attached to dissected myocardium | 72
source of embolism | 72
color flow Doppler interrogation | 72
diastolic flow in the apical cavity | 72
pulse wave Doppler | 72
diastolic flow into the apical cavity and systolic flow out of it | 72
cyclophosphamide therapy | 72
partial response | 72
reduction of the eosinophil count | 72
hypereosinophilic syndrome | 72
hypereosinophilia | 72
organ damage or dysfunction | 72
HES due to T-cell lymphoma | 72
cardiac complications of HES | 72
acute necrotic stage | 72
thrombotic stage | 72
fibrotic stage | 72
EM presents in stage 1 | 72
chest pain | 72
mimicking an acute myocardial infarction | 72
electrocardiogram | 72
ST-segment changes of ischemia | 72
embolic brain event | 72
intracardiac thrombus | 72
advances in echocardiography | 72
higher level of sensitivity | 72
cardiac masses | 72
differentiation between EM and apical mural thrombus | 72
CMR yields a respective sensitivity and specificity | 72
EM is typically characterized | 72
extensive myocardial hyperintensity on T2-weighted imaging | 72
subendocardial late enhancement | 72
endomyocardial biopsy | 72
gold standard for the diagnosis of EM | 72
partial or complete response | 72
corticosteroids | 72
monotherapy | 72
palliation | 72
multidisciplinary team meeting | 72
deterioration and poor prognosis | 72