12 years old | 0
male | 0
admitted to the hospital | 0
trauma to right ankle | -72
pain | -72
swelling of right ankle | -72
cough | -120
fever | -120
febrile | 0
tachycardia | 0
respiratory rate 25/min | 0
mildly swollen right ankle | 0
redness | 0
local rise of temperature | 0
tenderness over lateral malleolus | 0
restriction of ankle movements | 0
no neurovascular deficits | 0
plain X-ray of right ankle with leg normal | 0
haemoglobin-12.5gm% | 0
total count- 21.28K/uL | 0
neutrophils-19.77K/uL | 0
lymphocytes-0.75K/uL% | 0
CRP- 360.1mg/L | 0
ESR--60mm/hr | 0
RAfactor-negative | 0
ASO-titre- 400IU/ML | 0
sickling-negative | 0
urine routine normal | 0
admitted for treatment of suspected cellulitis | 0
pediatric opinion sought for cough | 0
Chest X-ray revealed pneumonia | 0
started on IV Cloxacillin 1gm four times daily | 0
blood culture revealed growth of Staphylococcus aureus | 24
sensitive to Cloxaciilin | 24
general condition deteriorated | 72
persistently elevated temperature | 72
tachycardia | 72
respiratory rate at 40/min | 72
SPO2- 87% at room air | 72
moderate swelling on whole of right leg | 72
tender calf | 72
positive Homan sign | 72
D-Dimer test negative | 72
CT angiogram of chest carried out | 72
no evidence of embolism | 72
right sided pleural effusion | 72
bilateral patchy pneumonia | 72
duplex scan of right lower limb suggestive of popliteal vein thrombosis | 72
thrombophilia work up for protein C &S | 72
anti-thrombin III negative | 72
treated with low molecular heparin | 72
treated with IV cloxacillin | 72
improved clinically | 120
calf swelling reduced | 120
blood parameters reverting to normalcy | 120
discharged | 336
treated with warfarin | 336
repeat duplex scan at 6 weeks normal | 504
followed up for period of 6 months | 1008
no signs of recurrence | 1008