84 years old | 0
woman | 0
chronic kidney disease | 0
hypertension | 0
mild cognitive dysfunction | 0
uterine mass | 0
presented to a regional hospital | -48
fever | -48
dry cough | -48
dyspnea | -48
chest x-ray | 0
bilateral lower lung patches | 0
pleural effusion | 0
septic shock | 0
acute kidney injury | 0
respiratory failure | 0
antibiotics | 0
fluid resuscitation | 0
tracheal intubation | 0
transferred to a tertiary hospital | 0
admitted to the intensive care unit | 0
curved gram-negative bacteria isolated from blood culture | 0
direct gram stain of pleural fluid | 0
curved gram-negative bacilli | 0
biochemical phenotype oxidase-positive | 0
catalase-negative | 0
urease-negative | 0
glucose-nonfermenting | 0
VITEK MS failed to identify | 0
VITEK2 GN ID card reported Burkholderia mallei | 0
16S rRNA PCR assay | 0
primers 11F | 0
primers 1512R | 0
amplified 16S rRNA genes | 0
1.5-kb amplified fragments from blood culture | 0
1.5-kb amplified fragments from pleural effusion culture | 0
identified as Paludibacterium purpuratum | 0
99.3% similarity | 0
98.9% similarity | 0
pleural effusion culture did not yield any bacteria | 0
16S rRNA sequencing identified P. purpuratum | 0
pneumonia | 0
empyema | 0
ampicillin-sulbactam | 0
bilateral pleural drainage | 0
24-Fr chest tubes | 0
extubated | 96
acute kidney injury resolved | 96
discharged home | 480
analyses of 16S rRNA sequences | 0
P. purpuratum strain B53371 | 0
99.6% similarity with P. purpuratum KJ031 | 0
98.3% similarity with P. yongneupense NBRC 106427 | 0
98.2% similarity with P. paludis KBP-21 | 0
whole-genome sequencing | 0
PaciBio Sequencing Platform | 0
genome size 3.63 M | 0
morphology assay | 0
drug susceptibility assay | 0
metabolic abilities assay | 0
grow on blood agar plate | 0
grow on chocolate agar plates | 0
gram stain showed curved gram-negative bacilli | 0
indole test negative | 0
hanging drop motility test negative | 0
growth less at 42°C | 0
no growth on MacConkey plate | 0
no growth on colistin nalidixic acid blood agar plate | 0
colony morphology on blood agar plate | 0
colony morphology on chocolate agar plate | 0
low MIC levels for ampicillin/sulbactam | 0
low MIC levels for piperacillin/tazobactam | 0
low MIC levels for cefotaxime | 0
low MIC levels for cefepime | 0
low MIC levels for fluoroquinolones | 0
low MIC levels for meropenem | 0
low MIC levels for aminoglycosides | 0
high MIC level for colistin | 0
phenotype microarray plates | 0
metabolize carbon sources | 0
metabolize nitrogen sources | 0
metabolize phosphorus sources | 0
metabolize sulfur sources | 0
utilize 33 substrates | 0
infection through inhalation | 0
misidentified by VITEK2 GN ID card | 0
Burkholderia mallei probability 90% | 0
ICR-Mo colistin resistance | 0
recovery with ampicillin/sulbactam therapy | 0
first invasive P. purpuratum infection in Taiwan | 0
exposure or inhalation of pathogen | 0
hypertension |;0
