60 years old| 0
    male|0
    emphysematous pyelonephritis|0
    diabetes mellitus|0
    failed renal allograft|0
    maintenance hemodialysis|0
    fever|0
    diffuse abdominal pain|0
    elevated white blood cell count|0
    computed tomographic scan showing air in failed renal allograft|0
    focal segmental glomerulosclerosis|- (prior to admission, exact time not specified)
    end-stage renal disease in 1990s|- (prior to admission, exact time not specified)
    dilated cardiomyopathy in mid-1990s|- (prior to admission, exact time not specified)
    bilateral radical nephrectomies for kidney cancer (right side in 1997, left in 1999)|- (prior to admission, exact time not specified)
    deceased donor renal transplant in 2001|- (prior to admission, exact time not specified)
    worsening left ventricular function in 2001|- (prior to admission, exact time not specified)
    ejection fraction of 25%|- (prior to admission, exact time not specified)
    severe mitral regurgitation|- (prior to admission, exact time not specified)
    acute renal failure in 2004|- (prior to admission, exact time not specified)
    transplant ureteric stricture in 2004|- (prior to admission, exact time not specified)
    balloon dilatation in 2004|- (prior to admission, exact time not specified)
    stent insertion in 2004|- (prior to admission, exact time not specified)
    transplant ureterectomy in 2004|- (prior to admission, exact time not specified)
    pyelovesicostomy of allograft in 2004|- (prior to admission, exact time not specified)
    psoas hitch of the bladder in 2004|- (prior to admission, exact time not specified)
    myocardial infarction in 2009|- (prior to admission, exact time not specified)
    medical therapy without revascularization in 2009|- (prior to admission, exact time not specified)
    transplant failure|- (prior to admission, exact time not specified)
    anuria|- (prior to admission, exact time not specified)
    hemodialysis|- (prior to admission, exact time not specified)
    deceased donor transplant wait list|- (prior to admission, exact time not specified)
    admission to ICU in 2012|- (prior to admission, exact time not specified)
    hypoglycemia in 2012|- (prior to admission, exact time not specified)
    fever in 2012|- (prior to admission, exact time not specified)
    non-ST-elevation myocardial infarction in 2012|- (prior to admission, exact time not specified)
    in-hospital arrest in 2012|- (prior to admission, exact time not specified)
    hepatomegaly in 2012|- (prior to admission, exact time not specified)
    elevated white blood cell count in 2012|- (prior to admission, exact time not specified)
    blood culture grew Bacteroides in 2012|- (prior to admission, exact time not specified)
    ciprofloxacin treatment|- (prior to admission, exact time not specified)
    metronidazole treatment|- (prior to admission, exact time not specified)
    CT scan of abdomen and pelvis|- (prior to admission, exact time not specified)
    piperacillin-tazobactam treatment|- (prior to admission, exact time not specified)
    transfer to tertiary care center|0
    hemodynamic stabilization|0
    emergent subcapsular nephrectomy|0
    necrotic kidney with pus encountered|0
    no significant blood loss|0
    postoperative transfer to ICU|0
    stable postoperatively|0
    death on postoperative day 4|96
    myocardial infarction on postoperative day 4|96
    histopathology showing necrotic kidney with acute inflammation|96
    total effacement of kidney architecture|96
    <|eot_id|>
    