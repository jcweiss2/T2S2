40 years old | 0
male | 0
admitted to the hospital (ICU) | 0
sepsis | 0
immunocompromised | 0
poorly controlled diabetes mellitus | 0
right thigh cellulitis | 0
diabetic ketoacidosis (DKA) | 0
developed inferior wall myocardial infarction | 0
developed right ventricular dysfunction | 0
altered sensorium | 0
hemodynamically unstable | 0
respiratory distress | 0
management of DKA | 0
management of acute coronary syndrome | 0
dual anti-platelets | 0
heparin | 0
statins | 0
invasive mechanical ventilation | 0
central line placement | 0
IV fluid resuscitation | 0
guided by two-dimensional echocardiography | 0
lung ultrasonography | 0
hemodynamic parameters | 0
oxygenation parameters | 0
vasoactive drugs | 0
anti-platelets | 0
therapeutic heparinization | 0
IV insulin infusion for glycemic control | 0
emphasis on electrolytes | 0
prolonged ICU stay | 0
neuromuscular weakness | 0
nosocomial infections | 0
ischemic cardiomyopathy | 0
developed grade III sacral bedsore | 0
Sphingobacterium multivorum bacteremia | 1008
cultured from peripheral blood | 1008
episode of high-grade fever | 1008
probable source (grade IV infected sacral bedsore) | 1008
sensitivity to piperacillin/tazobactam | 1008
sensitivity to levofloxacin | 1008
resistant to ceftazidime | 1008
resistant to amikacin | 1008
resistant to imipenem | 1008
resistant to carbapenem | 1008
resistant to aztreonam | 1008
treated with TMP/SMX | 1008
sensitive to TMP/SMX | 1008
diabetic ketoacidosis (DKA) |0
developed right ventricular dysfunction |0
altered sensorium |0
hemodynamically unstable |0
respiratory distress |0
management of DKA |0
management of acute coronary syndrome |0
dual anti-platelets |0
heparin |0
statins |0
invasive mechanical ventilation |0
central line placement |0
IV fluid resuscitation |0
guided by two-dimensional echocardiography |0
lung ultrasonography |0
hemodynamic parameters |0
oxygenation parameters |0
vasoactive drugs |0
anti-platelets |0
therapeutic heparinization |0
IV insulin infusion for glycemic control |0
emphasis on electrolytes |0
prolonged ICU stay |0
neuromuscular weakness |0
nosocomial infections |0
ischemic cardiomyopathy |0
developed grade III sacral bedsore |0
Sphingobacterium multivorum bacteremia |1008
cultured from peripheral blood |1008
episode of high-grade fever |1008
probable source (grade IV infected sacral bedsore) |1008
sensitivity to piperacillin/tazobactam |1008
sensitivity to levofloxacin |1008
resistant to ceftazidime |1008
resistant to amikacin |1008
resistant to imipenem |1008
resistant to carbapenem |1008
resistant to aztreonam |1008
treated with TMP/SMX |1008
sensitive to TMP/SMX |1008
