73 years old | 0
male | 0
admitted to the hospital | 0
jaundice | -72
2-cm mass in the pancreas | -72
obstruction of the common bile duct | -72
obstruction of the pancreatic duct | -72
no signs of metastases | -72
endoprosthesis placed endoscopically | -72
brush cytology | -72
adenocarcinoma | -72
severe progressive muscle weakness | -24
muscle weakness of legs | -24
muscle weakness of arms | -24
no pain | -24
no loss of sensation | -24
no skin abnormalities | -24
confined to a wheelchair | -24
diabetes mellitus type 2 | -672
spontaneous subdural hematoma | -672
surgically drained | -672
breast carcinoma in parents | -10000
colon carcinoma in parents | -10000
creatinine kinase level 12,570 U/l | 0
aspartate aminotransferase 594 U/l | 0
alanine aminotransferase 523 U/l | 0
lactate dehydrogenase 648 U/l | 0
C-reactive protein 11 mg/l | 0
magnetic resonance imaging | 0
diffuse edema in upper leg muscles | 0
diffuse edema in lower leg muscles | 0
inflammatory process | 0
muscle biopsy | 0
necrotic fibers | 0
macrophages | 0
regenerating fibers | 0
membrane attack complex positive fibers | 0
MHC-I positive non-necrotic muscle fiber | 0
skin histology | 0
no skin abnormalities | 0
dexamethasone therapy | 0
prednisone therapy | 0
intravenous immunoglobulin | 0
laparoscopic pancreatoduodenectomy | 10
R0 resected pT3N0M0 distal cholangiocarcinoma | 10
no adjuvant chemotherapy | 10
improvement in NAM symptoms | 24
muscle strength increased | 24
able to walk a few steps | 38
pancreatic fistula | 10
percutaneous drain | 10
pneumonia | 42
treated with antibiotics | 42
deteriorated general condition | 42
confined to a wheelchair | 42
admitted to intensive care unit | 84
pneumosepsis | 84
maximized supportive care | 84
enteral tube feeding | 84
no signs of recovery | 112
discontinuation of medical treatment | 112
death | 128