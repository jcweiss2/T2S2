23 years old | 0
postpartum woman | 0
septic shock | 0
admitted to the intensive care unit | 0
severe iron deficiency anemia | -672
gestational hypertension | -672
meconium-stained amniotic fluid | -672
prolonged rupture of the membranes | -672
chorioamnionitis | -48
urgent cesarean section | -48
purulent postpartum endometritis | -24
fever | -24
chills | -24
purulent uterine discharge | -24
fundal tenderness | -24
arterial line placement | -24
blood culture | -24
sepsis | -12
septic shock | -12
organ failure | -12
SOFA score 16-20 | -12
ARDS | -12
acute respiratory distress syndrome | -12
norepinephrine infusion | -12
dobutamine infusion | -6
left ventricular systolic dysfunction | -6
ejection fraction 32% | -6
mottled fingers and toes | -6
mottled abdominal wall | -6
hysterectomy | -48
transfer to hospital | 0
massive aseptic necrosis of fingers | 0
massive aseptic necrosis of toes | 0
massive aseptic necrosis of metatarsal region | 0
massive aseptic necrosis of anterior abdominal wall | 0
sepsis-induced multiple system failure | 0
ARDS | 0
encephalopathy | 0
systolic heart failure | 0
acute kidney injury | 0
invasive blood pressure 100/70 mmHg | 0
heart rate 150/min | 0
arterial oxygen saturation 85-92% | 0
body temperature 38.4°C | 0
sedation with dexmedetomidine | 0
mechanical ventilation | 0
crackles over the right middle and lower zones of the lungs | 0
hemodynamic support with norepinephrine | 0
hemodynamic support with dobutamine | 0
Hb 9 g/dl | 0
WBC 22 × 10^9/L | 0
C-reactive protein 200.5 mg/L | 0
lactate 4 mmol/L | 0
procalcitonin 32 ng/ml | 0
сreatine-kinase MB 15.1 IU/L | 0
BNP 5,000 ng/ml | 0
platelets 90 × 10^9/L | 0
fibrinogen 114 mg/dl | 0
activated partial thromboplastin time 128 s | 0
international normalized ratio 1.27 | 0
prothrombin time 16.9 s | 0
transthoracic echocardiography | 0
reduced ejection fraction 38% | 0
bilateral infiltrations on chest radiography | 0
mild acute respiratory distress syndrome | 0
PaO2/FiO2 250 mmHg | 0
blood culture with multiple drug-resistant Escherichia coli | 0
blood culture with Pseudomonas aeruginosa | 0
blood culture with Acinetobacter baumannii | 0
antibacterial therapy | 0
goal-directed fluid therapy | 0
nutritional support | 0
protective mechanical ventilation | 0
hydrocortisone | 0
fresh frozen plasma | 0
high dose of ascorbic acid and thiamine | 0
skin wound management with dressing and moist healing products | 0
weaning off mechanical ventilation | 168
weaning off vasopressor therapy | 168
no neurological consequences | 168
end-organ functions returned to normal | 168
necrotic masses debrided | 240
autodermoplasty | 240