79 years old | 0
male | 0
Chinese ethnicity | 0
COPD | 0
stable ischaemic heart disease | 0
bicytopenia | -168
normocytic, normochromic anemia | -168
decreased reticulocyte response | -168
leukopenia | -168
bone marrow aspirate | -168
mild dysplastic changes | -168
plasmacytosis | -168
bone marrow trephine | -168
increased number of CD 138+ plasma cells | -168
hernia repair | -168
admitted to the hospital | 0
dyspnoea | 720
fever | 720
anemic | 720
leukopenic | 720
treated for possible neutropenic sepsis | 720
pneumonia | 720
mild congestive cardiac failure | 720
acute infective exacerbation of COPD | 720
cultures from blood, urine, stool, and sputum | 720
TB PCR and AFB smears | 720
chest X-ray | 720
small bilateral pleural effusions | 720
focal consolidation in bilateral midzones | 720
carbapenem antibiotic | 720
transfusion support | 720
serum electrophoresis and immunofixation | 720
no conclusive evidence of a monoclonal paraprotein | 720
faint bands at IgM and lambda lanes | 720
urine IFE at lambda lane | 720
serum M-band | 720
skeletal survey | 720
serum calcium | 720
flow cytometry of peripheral blood | 720
polyclonal, circulating lymphoplasmacytoid cells | 720
CT scan of neck/chest/abdomen/pelvis | 720
mild splenomegaly | 720
small volume lymphadenopathy | 720
HIV serology | 720
negative | 720
repeat bone marrow studies | 720
deferred | 720
developed another fever | 744
broad-spectrum antimicrobials | 744
chest X-ray | 744
bilateral pleural effusions | 744
pleurocentesis | 744
bloody pleural fluid | 744
bronchoscopic evaluation | 744
connective tissue disease workup | 744
unremarkable | 744
BAL studies | 744
negative for malignancy and tuberculosis | 744
atypical plasma cells | 744
fungal elements | 744
morphology of a mixture of Candida and Cryptococcus | 744
serum cryptococcal antigen | 744
negative | 744
hypotensive | 744
admitted to the Intensive Care Unit | 744
inotropic support | 744
GCSF | 744
intravenous Amphotericin B | 744
presumptive diagnosis of disseminated cryptococcosis | 744
Amphotericin | 744
changed to IV Ambisome | 768
worsening renal function | 768
pericardial effusion | 768
stable | 768
cryptococcal involvement | 768
pericardiocentesis | 768
deferred | 768
BAL cultures | 768
grew CN | 768
sensitive to fluconazole | 768
Ambisome | 768
changed to IV Fluconazole | 768
deteriorated | 816
passed away | 816
bone marrow biopsy specimen | 816
reexamined | 816
GMS stain | 816
revealed two large cells containing GMS-positive yeast-like structures | 816
identical to those detected in BAL | 816
confirmed to be CN via PCR | 816
diagnosis of chronic disseminated CN infection | 816
pleural and pericardial effusion | 816
lymph node | 816
lung | 816
bone marrow involvement | 816