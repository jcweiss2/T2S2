61 years old | 0
African American female | 0
admitted to the hospital | 0
end-stage renal disease | -6720
adult polycystic kidney disease | -6720
living-related kidney transplant | -6720
fever | -120
gastrointestinal symptoms | -120
diarrhea | -120
nausea | -120
attended a funeral | -240
hypertension | 0
gout | 0
histoplasmosis | 0
tacrolimus | -6720
mycophenolate mofetil (MMF) | -6720
prednisone | -6720
itraconazole | -6720
allopurinol | -6720
labetalol | -6720
hydralazine | -6720
febrile | 0
pulse rate 87 beats per minute | 0
blood pressure 151/85 mm Hg | 0
respiratory rate 24 breaths per minute | 0
oxygen saturation 92% to 97% on room air | 0
respiratory distress | 0
decreased breath sounds on the left side of the chest | 0
mild mid to lower lung infiltrate bilaterally | 0
mild mid to lower lung infiltrate on the left side | 0
mild mid to lower lung infiltrate on the right side | 0
few scattered rounded ground glass and consolidative opacities | 0
segmental lung consolidation | 0
COVID-19 testing positive | 0
ceftriaxone | 0
azithromycin | 0
intravenous fluids | 0
antipyretics | 0
MMF held | 0
tacrolimus continued | 0
prednisone continued | 0
oxygen therapy | 0
fever resolved | 24
discharged | 120
MMF restarted | 120 
immunosuppressive regimen continued | 120 
doing well | 336