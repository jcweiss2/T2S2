40 years old | 0
female | 0
obesity | 0
confusion | -168
dysuria | -168
left EPN | -168
CT scan | -168
admitted to Medical Intensive Care Unit (ICU) | 0
awake and oriented | 0
denied hematuria | 0
denied flank pain | 0
denied chest pain | 0
denied shortness of breath | 0
denied history of nephrolithiasis | 0
afebrile | 0
tachycardic | 0
normotensive | 0
tachypneic | 0
saturating well on room air | 0
WBC of 34 | 0
platelet count 66 | 0
lactate 5.8 | 0
BUN 56 | 0
creatinine 3.22 | 0
glucose 485 | 0
alkaline phosphatase 498 | 0
AST 39 | 0
ALT 43 | 0
Hemoglobin A1C 7.6 | 0
urine and blood cultures grew E. coli | 0
suprapubic tenderness | 0
gas within the parenchyma of the upper left kidney | 0
4 mm stone within the proximal left ureter | 0
air in the collecting systems of both kidneys | 0
heterogenous liver with cirrhotic nodules | 0
moderate amount of abdominal ascites | 0
diagnosed with Child Class C cirrhosis | 0
started on rifaximin and lactulose | 0
nonalcoholic fatty liver disease | 0
Model for End-Stage Liver Disease (MELD-Na) score 31 | 0
guarded prognosis | 0
intravenous fluids | 0
insulin drip | 0
Zosyn | 0
insertion of bilateral double J stents | 12
retrograde pyelogram | 12
no evidence of hydroureteronephrosis | 12
foley left in place | 12
worsening acidosis | 24
required continued intubation | 24
required dialysis | 72
required bicarbonate drip | 72
required pressors | 72
tachypnea | 72
low volumes | 72
repeat CT scan | 72
worsening left EPN | 72
near complete necrosis of the left renal upper pole | 72
new right EPN | 72
new right colon pneumatosis | 72
portal venous gas | 72
planning for definitive surgical intervention | 72
emergent left nephrectomy | 72
general surgery consulted | 72
necessity of bowel resection | 72
comfort measures | 96
terminally extubated | 96
died | 96