31 years old | 0
male | 0
admitted to ICU | 0
postexploratory laparotomy | -72
right thoracotomy | -72
gunshot wound to the abdomen and chest | -72
left arm injury | -72
left elbow fracture | -72
open reduction internal fixation (ORIF) | -72
septic shock | -72
acute kidney injury | -72
chest infection | 0
infected laparotomy wound | 0
piperacillin/tazobactam therapy | 0
continuous fever | 0
leukocytosis | 0
persistent source of infection | 0
abdominal wound | 0
left-hand ORIF site wound | 0
frequent dressing and debridement | 0
P. stuartii isolates identified | 0
carbapenem-resistant P. stuartii isolate detected | 528
resistant to ciprofloxacin | 528
resistant to trimethoprim/sulfamethoxazole | 528
resistant to gentamicin | 528
resistant to imipenem | 528
resistant to meropenem | 528
sensitive to amikacin | 528
highly febrile | 720
piperacillin/tazobactam 4.5 g provided iv | 720
fever persistent | 744
leukocytes increasing | 744
septic screening | 744
piperacillin/tazobactam changed to meropenem | 744
growth of P. stuartii and carbapenem-resistant K. pneumoniae in urine | 840
growth of P. stuartii and carbapenem-resistant K. pneumoniae in wound | 840
growth of P. stuartii and carbapenem-resistant K. pneumoniae in blood | 840
tracheal aspirate culture report | 888
carbapenem-resistant P. stuartii isolate resistant to amikacin | 888
carbapenem-resistant P. stuartii isolate resistant to ciprofloxacin | 888
carbapenem-resistant P. stuartii isolate resistant to trimethoprim/sulfamethoxazole | 888
carbapenem-resistant P. stuartii isolate resistant to gentamicin | 888
carbapenem-resistant P. stuartii isolate intermediate to meropenem | 888
meropenem dosing regimen changed | 888
colistin prescribed | 888
follow-up septic screen | 1056
growth of multidrug-resistant Acinetobacter baumannii in left-hand ORIF site wound | 1128
growth of multidrug-resistant Acinetobacter baumannii in tracheal aspirate | 1128
chest X-ray ordered | 1128
meropenem and colistin discontinued | 1344
transferred to ward | 1344
stable with no signs and symptoms of infection | 1344