20 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
non-smoker | 0 | 0 | Factual
occupational smoke exposure | -336 | 0 | Factual
fever | -336 | 0 | Factual
productive cough | -336 | 0 | Factual
night sweats | -336 | 0 | Factual
malaise | -336 | 0 | Factual
myalgia | -336 | 0 | Factual
treated with roxithromycin | -168 | -24 | Factual
no clinical response | -24 | 0 | Factual
admitted to the hospital | 0 | 0 | Factual
temperature 38.4°C | 0 | 0 | Factual
blood pressure 130/70 mmHg | 0 | 0 | Factual
pulse 88 bpm | 0 | 0 | Factual
oxygen saturation 97% | 0 | 0 | Factual
dyspnoea | 0 | 0 | Factual
tachypnoea | 0 | 0 | Factual
bronchial breathing sounds | 0 | 0 | Factual
crackles over the right lung | 0 | 0 | Factual
white blood cells 11.54×10^3/μl | 0 | 0 | Factual
total eosinophils 92×10^4/μl | 0 | 0 | Factual
haemoglobin 13.7 g/dl | 0 | 0 | Factual
creatinine 1.1 mg/dl | 0 | 0 | Factual
C-reactive protein (CRP) 11 mg/dl | 0 | 0 | Factual
liver enzymes elevated | 0 | 0 | Factual
ALP 524 | 0 | 0 | Factual
GGT 320 | 0 | 0 | Factual
ALT 406 | 0 | 0 | Factual
AST 137 | 0 | 0 | Factual
abdominal ultrasound normal | 0 | 0 | Factual
chest radiograph showed infiltrates | 0 | 0 | Factual
treated with IV cefuroxime | 0 | 48 | Factual
blood and sputum cultures negative | 0 | 48 | Factual
urine Legionella antigen test negative | 0 | 48 | Factual
persistent high-grade fever | 48 | 96 | Factual
antibiotic treatment changed to moxifloxacin | 48 | 48 | Factual
respiratory distress | 96 | 120 | Factual
oxygen saturation dropped to 88% | 96 | 96 | Factual
arterial blood gas disclosed PaO2 67 mmHg | 96 | 96 | Factual
CRP increased to 14 mg/dl | 96 | 96 | Factual
liver enzymes elevated | 96 | 96 | Factual
leucocytosis 12.8×10^3/μl | 96 | 96 | Factual
eosinophil count 1.33×10^3 cells/μl | 96 | 96 | Factual
follow-up chest radiogram showed progression | 96 | 96 | Factual
diffuse bilateral infiltrates | 96 | 96 | Factual
intubated | 120 | 120 | Factual
mechanically ventilated | 120 | 120 | Factual
transferred to the intensive care unit | 120 | 120 | Factual
broncho-alveolar lavage demonstrated 30% eosinophils | 144 | 144 | Factual
diagnosed with AEP | 144 | 144 | Factual
IV glucocorticoids administered | 144 | 144 | Factual
prompt improvement | 144 | 168 | Factual
resolution of fever | 144 | 168 | Factual
successful extubation | 168 | 168 | Factual
chest radiogram showed regression of bilateral infiltrates | 168 | 168 | Factual
eosinophil count dropped to 260 cells/μl | 168 | 168 | Factual
discharged | 216 | 216 | Factual
oral prednisone 60 mg/day | 216 | 216 | Factual
tapering over 3 months | 216 | 744 | Factual