67 years old|0
woman|0
sternoclavicular septic arthritis|0
recurrent bacteremia|0
previous bacterial endocarditis|0
end-stage renal disease|0
hemodialysis|0
persistent cough|0
dysphagia to solid foods|0
large, true aneurysm of the proximal right subclavian artery|0
proximity to the clavicular infection|0
mSAA|0
cardiac clearance obtained|0
open repair|0
partial median sternotomy|0
right infraclavicular extension|0
partial right claviculectomy|0
clavicle reconstruction deferred|0
highly inflamed and fibrous mediastinal/periclavicular tissue|0
right internal jugular vein ligated and divided|0
multiple enlarged collateral veins ligated and divided|0
excision of the aneurysm|0
right phrenic nerve identified and protected|0
right vertebral artery identified|0
innominate-to-right subclavian arterial bypass|0
reimplantation of the right common carotid artery|0
rifampin-soaked, Dacron graft used|0
specimens sent for pathologic analysis|0
postoperative head and neck edema|0
endotracheal ventilation|0
extubated|168
transferred out of intensive care unit|216
discharged|480
chronic osteomyelitis of the clavicular head|0
partial wall necrosis|0
organized thrombus|0
methicillin-sensitive Staphylococcus aureus|0
6-week course of intravenous cefazolin|0
converted to cephalexin|0
free from recurrent bacteremia|0
no residual head or neck edema|0
minimal change in upper extremity functioning|0
denies vasculogenic symptoms|0
