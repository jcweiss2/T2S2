25 years old | 0 | 0 
female | 0 | 0 
housewife | 0 | 0 
admitted to the hospital | 0 | 0 
given birth | -24 | -24 
spontaneous vaginal delivery | -24 | -24 
episiotomy | -24 | -24 
severe pain | -24 | 0 
shortness of breath | -24 | 0 
worsening pain | -24 | 0 
tachypnea | 0 | 0 
oxygen saturation 56% | 0 | 0 
high-flow oxygen supply | 0 | 24 
tachycardia | 0 | 0 
pulse 121 bpm | 0 | 0 
afebrile | 0 | 0 
blood pressure unrecordable | 0 | 0 
hypotensive | 0 | 24 
noradrenaline infusion | 0 | 24 
IV heparin | 0 | 0 
IV amoxicillin-clavulanate | 0 | 0 
transferred to tertiary hospital | 0 | 0 
elective intubation | 0 | 0 
severe metabolic acidosis | 0 | 0 
lactic acidosis | 0 | 24 
worsening respiratory distress | 0 | 0 
crystalloid | 0 | 24 
inotropes | 0 | 24 
adrenaline | 0 | 24 
vasopressin | 0 | 24 
dobutamine | 0 | 24 
grossly swollen right thigh | 0 | 0 
extensive blistering ecchymotic patches | 0 | 0 
necrotizing fasciitis | 0 | 24 
septicemic shock | 0 | 24 
acute kidney injury | 0 | 24 
rhabdomyolysis | 0 | 24 
coagulopathy | 0 | 24 
thrombocytopenia | 0 | 24 
ischemic hepatitis | 0 | 24 
IV meropenem | 0 | 24 
IV clindamycin | 0 | 24 
IV vancomycin | 0 | 24 
high vaginal swab | 0 | 0 
CT pulmonary angiography | 0 | 0 
pulmonary embolism | 0 | 0 
bedside echocardiography | 0 | 0 
intravenous immunoglobulin | 0 | 120 
toxin neutralization | 0 | 120 
continuous veno-venous hemofiltration | 0 | 168 
lactate 9.8-18 mmol/L | 0 | 168 
creatinine kinase 29783 U/L | 0 | 168 
skin lesion spread | 24 | 168 
blistering of bilateral lower limbs | 24 | 168 
bluish discoloration | 24 | 168 
Gram positive cocci in chains | 24 | 24 
S. pyogenes | 24 | 24 
multidisciplinary discussion | 144 | 144 
group A streptococcal toxic shock syndrome | 144 | 168 
IV crystalline penicillin G | 144 | 168 
toxin suppression | 144 | 168 
surgical intervention | 168 | 168 
skin biopsy | 168 | 168 
death | 168 | 168 
septic shock | 168 | 168 
tissue necrosis | 168 | 168 
toxic shock syndrome | 168 | 168 
S. pyogenes | 168 | 168