70 years old | 0
    woman | 0
    presented to emergency | 0
    acute abdominal pain | 0
    immunocompromised | 0
    type II diabetes | 0
    previous splenectomy | -315360
    trauma | -315360
    multiple previous laparotomies | 0
    adhesive bowel obstruction | 0
    CT abdomen | 0
    perforated splenic flexure malignancy | 0
    laparotomy | 0
    grossly dilated large bowel | 0
    no obvious perforation | 0
    loop colostomy | 0
    decompression of large colon | 0
    intravenous Piperacillin/Tazobactam | 0
    vancomycin | 0
    fluconazole | 0
    admitted to intensive care unit | 0
    ongoing shock | 0
    high vasopressor requirement | 0
    noradrenaline requirement | 0
    erythematous patch on left thigh | 14
    creatine kinase of 19000 | 14
    bedside finger test | 14
    dirty dishwater fluid | 14
    necrotic fat | 14
    lack of bleeding | 14
    taken to theatre for urgent debridement | 14
    suspected NF | 14
    antibiotics changed to Meropenem | 14
    Vancomycin | 14
    Lincomycin | 14
    Fluconazole | 14
    extensive debridement of soft tissue on left thigh | 14
    muscle involvement | 14
    radiological evidence of disease progression | 24
    gas in muscle compartments on lower limb X-rays | 24
    CT abdomen and lower limbs demonstrating gas | 24
    non-contiguous area in right gluteal region | 24
    diagnosis of multi-focal non-contiguous necrotising myositis | 24
    multiple comorbidities | 24
    very high mortality risk | 24
    low risk of recovery | 24
    palliated | 24
    swab | 24
    tissue microscopy | 24
    no pathogen isolated | 24
    early commencement of broad-spectrum antibiotics | 0
    