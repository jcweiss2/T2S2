28 years old | 0
    male | 0
    admitted to the hospital | 0
    gingival swelling | 0
    AML [t(9;11)(p22;q23); MLLT3(AF9)-MLL] diagnosis | -21600
    bone marrow aspiration | -21600
    peripheral blood stem cell transplantation (PBSCT) | -16320
    HLA-identical sibling donor | -16320
    conditioning regimen (busulfan 12.8 mg/kg, cyclophosphamide 120 mg/kg) | -16320
    GVHD prophylaxis (cyclosporine A, short-term methotrexate) | -16320
    grade I acute GVHD | -16320
    methylprednisolone (1 mg/kg) | -16320
    cyclosporine A discontinuation | -12960
    molecular relapse of AML | -12960
    bridging therapies (azacitidine, gemtuzumab ozogamicin) | -12960
    donor lymphocyte infusion | -12960
    molecular complete remission | -12960
    second bone marrow transplantation | -10560
    HLA-identical unrelated donor | -10560
    conditioning regimen (cyclophosphamide 120 mg/kg, total body irradiation 1200 cGy) | -10560
    GVHD prophylaxis (tacrolimus, short-term methotrexate) | -10560
    skin and gut GVHD | -10560
    cytomegalovirus enterocolitis | -10560
    discharged after second HSCT | -10560
    bronchiolitis obliterans | -7200
    high-dose pulse methylprednisolone therapy | -7200
    mycophenolate mofetil | -7200
    hematological relapse of AML | -8760
    admitted for salvage chemotherapy | 0
    recurrent pneumonia | 0
    watery diarrhea | 0
    maculopapular skin rash | 0
    infiltrative shadow in left lung on CT | 0
    meropenem | 0
    vancomycin | 0
    salvage chemotherapy (mitoxantrone, etoposide, intermediate-dose cytarabine) | 96
    diarrhea worsened | 240
    maculopapular skin rash expansion | 240
    intestinal edema on CT | 240
    white blood cells 20 /μL | 240
    hemoglobin 8.4 g/dL | 240
    platelets 12,000/μL | 240
    lactate dehydrogenase 228 U/L | 240
    C-reactive protein 1.24 mg/dL | 240
    Clostridium difficile toxins A/B negative | 240
    glutamate dehydrogenase (GDH) negative | 240
    suspected recurrence of acute gut GVHD | 240
    methylprednisolone increased to 120 mg/day | 240
    beclomethasone dipropionate 8 mg/day | 240
    diarrhea worsened | 312
    steroid pulse therapy (methylprednisolone 1 g/day for 3 days) | 312
    colonoscopy not possible | 312
    hemorrhagic diarrhea | 384
    blood cultures positive for Gram-negative bacilli | 384
    minocycline | 384
    ciprofloxacin | 384
    S. maltophilia identification | 408
    trimethoprim-sulfamethoxazole | 408
    died | 432
    respiratory failure progression | 432
    hemodynamic instability | 432
    hemorrhagic enterocolitis | 432
    pneumonia with septic shock | 432
    erosion in terminal ileum | 432
    petechial hemorrhaging in lower intestinal tract | 432
    Gram-negative bacilli in ileum layers | 432
    no apoptotic bodies | 432
    no CMV-infected cells | 432
    no pseudomembranous colitis | 432
    hemorrhagic pneumonia in left lung | 432
    no Gram-negative bacilli proliferation in other organs | 432
    

