68 years old | 0
man | 0
presented to the hospital | 0
subjective fever | 0
bilateral leg pain | 0
worsening blistering | 0
bleeding from BP lesions of the lower extremities | 0
chronic history of BP | -35040
BP diagnosed | -35040
hospital admission 2 weeks prior | -336
severe flare of BP | -336
prednisone 60 mg PO daily | -336
prolonged 6-week taper | -336
doxycycline 100 mg PO twice daily | -336
shave biopsy of the bullous skin lesions | -336
refractory CLL | 0
recurrent deep vein thrombosis | 0
apixaban 5 mg twice daily | 0
chronic obstructive pulmonary disease | 0
diastolic heart failure | 0
non-insulin dependent diabetes mellitus | 0
hypogammaglobulinemia | 0
intravenous immunoglobulin 400 mg/kg | 0
11q deletion CLL | -218400
treatment with R-CVP | -218400
treatment with FR | -218400
ibrutinib 420 mg PO daily | -26208
maintained on ibrutinib for approximately 3 years | -26208
initial vital signs were normal | 0
multiple round hyperpigmented macules on the trunk, upper and proximal lower extremities | 0
numerous necrotic ulcers with hemorrhagic keratotic eschars | 0
surrounding bullae from recent BP flare | 0
comprehensive metabolic profile within normal limits | 0
white blood cell count 2,600/µL | 0
absolute neutrophil count 1,100/µL | 0
hemoglobin 9.3 g/dL |1| 0
platelets 103,000/µL | 0
given intravenous immunoglobulin | 0
IgG of 350 mg/dL | 0
developed sepsis | 0
atrial fibrillation with rapid ventricular response | 0
hypotension | 0
transferred to the intensive care unit | 0
started on vancomycin 15 mg/kg intravenous every 12 h | 0
meropenem 1 g intravenous every 8 h | 0
ibrutinib held | 0
prophylactic acyclovir 400 mg PO twice daily continued | 0
prednisone tapered down to 20 mg PO daily | 0
shave biopsy results returned as trophozoites with concern for possible fungal infection | 0
started intravenous fluconazole 400 mg daily | 0
stabilized in the intensive care unit over several days | 0
atrial fibrillation controlled with metoprolol | 0
vancomycin discontinued | 0
meropenem discontinued | 0
new necrotic lesions continued to develop | 0
repeat punch biopsies performed | 0
switched to intravenous liposomal amphotericin B 5 mg/kg daily | 0
blood cultures negative | 0
cryptococcal antigen negative | 0
urine histoplasma antigen negative | 0
urine blastomycosis antigen negative | 0
serum coccidioides antibody negative | 0
computed tomography of the chest, abdomen and pelvis with contrast significant for hiatal hernia | 0
splenomegaly | 0
transferred out of the intensive care unit | 0
continued on intravenous liposomal amphotericin B | 0
appropriate wound care | 0
pain control | 0
punch biopsies showed septate hyphae with chains of arthroconidia | 0
x-rays of bilateral tibia and fibula unremarkable | 0
subcutaneous skin thickening consistent with BP | 0
fungal cultures from punch biopsies returned positive for mucormycosis | 336
extensive necrotic lesions with thick black eschars | 336
several lesions loosening and sloughing off | 336
bilateral magnetic resonance images negative for osteomyelitis | 336
no evidence of extension of mucormycosis beyond subcutaneous tissues | 336
plastic surgery consulted for debridement | 336
decision to continue with antifungal therapy and aggressive wound care | 336
developed foul smelling drainage with green tinge | 480
white blood cell count increased to 17,600/µL | 480
wound culture collected | 480
started on daptomycin 6 mg/kg daily | 480
meropenem 1 g every 8 h | 480
completed 7-day course with improvement | 480
wound cultures grew Pseudomonas | 480
wound cultures grew E. coli | 480
repeat blood cultures negative | 480
received 4 weeks of intravenous liposomal amphotericin B | 672
transitioned to posaconazole 400 mg PO twice daily | 672
wounds continued to gradually heal | 672
discharged to skilled nursing facility | 1344
