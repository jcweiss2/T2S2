73 years old | 0
male | 0
admitted to the hospital | 0
COVID-19 | -24
hypertension | -8760
diabetes mellitus | -8760
percutaneous coronary intervention (PCI) | -8760
aspirin | -8760
fever | -24
cough | -24
chest radiography | 0
ill-defined, hazy, and streaky density in both the lungs | 0
hydroxychloroquine treatment | 0
pneumonia | 0
hypotension | 24
melena | 24
tachycardia | 24
peripheral oxygen saturation (SpO2) of approximately 80% | 24
hemoglobin level had decreased to 6.3 mg/dl | 24
blood transfusion | 24
endotracheal intubation | 24
arterial catheter insertion | 24
central venous catheter insertion | 24
esophagogastroduodenoscopy (EGD) | 49
duodenal ulcer | 49
endoscopic hemoclipping and embolization | 73
abdominal pain | 97
subphrenic free air | 97
pneumoperitoneum | 97
exploratory laparotomy | 105
general anesthesia | 105
intubation | 105
mechanical ventilation | 105
invasive arterial blood pressure (ABP) monitoring | 105
electrocardiography (ECG) monitoring | 105
heart rate monitoring | 105
SpO2 monitoring | 105
bispectral index monitoring | 105
propofol | 105
rocuronium | 105
sevoflurane | 105
remifentanil | 105
lung-protective mechanical ventilation strategy | 105
surgery | 105
pyloric exclusion | 105
primary closure of the perforation | 105
gastrojejunostomy | 105
midazolam | 125
rocuronium | 125
transfer to the ward | 125
infection control | 125
disinfection | 125
sterilization | 125
septic shock | 153
norepinephrine | 153
expired | 168
SARS-CoV-2 | -24
RT-PCR | -24
nasopharyngeal and oropharyngeal swabs | 49
RT-PCR | 49
SARS-CoV-2 | 49
pneumonia | 49
C-reactive protein | 49
fever | 49
elevated C-reactive protein | 121
fever | 121
pneumonic infiltration | 121
pleural effusion | 121
septic shock | 153
hypotension | 153
norepinephrine | 153
expired | 168