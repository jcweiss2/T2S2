59 years old | 0
    male | 0
    admitted to the hospital | 0
    intermittent diarrhea | -120
    developed soon after eating contaminated food | -120
    reduced urine volume | -72
    diarrhea with water-like stools more than 10 times/d | -120
    abdominal pain | -120
    nausea | -120
    vomiting | -120
    decreased production of dark-colored urine (50-100 mL/d) | -72
    fatigue | -72
    limb weakness | -72
    transferred to the ICU | -72
    temperature 38.5 °C | 0
    pulse 128 beats/min | 0
    respiration 22 breaths/min | 0
    blood pressure 70/40 mmHg | 0
    no lung abnormalities | 0
    no cardiac abnormalities | 0
    slightly puffy abdomen | 0
    soft abdomen | 0
    upper abdominal pressure | 0
    back pain | 0
    bowel “chirping” 5-6 times/min | 0
    hemoglobin 18.3 g/dL | 0
    white blood cell count 21.4 × 10^9/L | 0
    71.9% neutral granulocytes | 0
    platelet count 169 × 10^9/L | 0
    metabolic acidosis | 0
    blood gas pH 7.35 | 0
    PCO2 30 mmHg | 0
    PO2 66 mmHg (FiO2 60%) | 0
    PO2/FiO2 110 mmHg | 0
    bicarbonate 16.6 mmol/L | 0
    base excess -9.0 mmol/L | 0
    lactate 3.5 mmol/L |    0
    aspartate aminotransferase 573.1 U/L | 0
    alanine aminotransferase 47 U/L | 0
    total bilirubin 7.58 µmol/L | 0
    serum creatinine 708.8 µmol/L | 0
    urea 20.48 mmol/L | 0
    albumin 26.9 g/L | 0
    prothrombin time 12.5 s | 0
    activated partial thromboplastin time 31.3 s | 0
    international normalized ratio 1.08 | 0
    procalcitonin 32.60 ng/mL | 0
    negative hepatitis tests (HBsAg, HBsAb, HBeAg, HBeAb, HBcAb, HCV) | 0
    negative autoimmune hepatitis tests (antinuclear antibodies, smooth muscle antigen, soluble liver antigen antibodies, liver-kidney microsome-1, other autoantibodies) | 0
    Salmonella not detected in stool culture | 0
    Shigella not detected in stool culture | 0
    Clostridium difficile toxin A toxin B negative | 0
    Gram-negative bacilli in stool | 0
    Gram-positive cocci in stool | 0
    empirical meropenem treatment | 0
    blood culture Klebsiella pneumoniae sensitive to meropenem | 0
    Klebsiella pneumoniae bacteraemia | 0
    sepsis | 0
    septic shock | 0
    acute kidney injury | 0
    APACHE II score 18 | 0
    SOFA score 10 | 0
    intravenous crystalloid fluid 2500 mL within first 3 h | 0
    invasive dynamic hemodynamic monitoring | 0
    blood pressure increased to 80/55 mmHg | 3
    noradrenaline administration | 3
    mean arterial pressure 65 mmHg | 3
    CRRT with oXiris® hemofilter | 0
    CVVHDF mode | 0
    12-French double-lumen catheter in right femoral vein | 0
    pre-dilution prescription | 0
    blood flow rate 150 L/min | 0
    regional citrate anticoagulation | 0
    mild hypocalcemia | 0
    intravenous calcium supplementation | 0
    meropenem continued | 0
    CRRT with oXiris® filter for 72 h | 72
    vital signs stable | 72
    infection well controlled | 72
    noradrenaline infusion reduced to 0.05 µg/kg per minute | 65
    noradrenaline stopped at 65 h | 65
    lactate level 2.1 mmol/L | 6
    lactate clearance rate 40% | 6
    endotoxin levels declined | 6
    IL-6 levels declined | 6
    IL-10 levels declined | 6
    PCT decreased to 4.98 ng/mL | 72
    urine volume gradually increased over 10 d | 240
    SCr decreased from 708.8 µmol/L to 241 µmol/L over 3 d | 72
    SOFA score decreased from 10 to 3 | 72
    APACHE II score decreased from 18 to 6 | 72
    hemodynamically stable | 72
    traditional filter (AN69 hemofilter) | 72
    intermittent CVVHDF | 72
    CRRT discontinued after kidney function recovery | 480
    significant amelioration of septic shock | 600
    discharged | 600
    kidney function returned to normal | 600
    