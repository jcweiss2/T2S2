61 years old | 0
male | 0
admitted to the hospital | 0
intermittent high-grade fever | -720
swelling of right knee joint | -720
severe pain | -720
inability to weight bear | -720
inability to walk due to knee pain | -168
treated for right knee pain | -720
treated for urinary tract infection | -720
type II diabetes mellitus | 0
sudden onset breathlessness | -24
conscious | 0
febrile | 0
tachycardic | 0
tachypnoeic | 0
hypotensive | 0
reduced saturation | 0
extensive bilateral crepitations | 0
right knee swelling | 0
warm | 0
tender | 0
septic arthritis right knee | 0
severe septicemia | 0
septic shock | 0
intubated | 0
fluid resuscitated | 0
inotropes | 0
vasopressors | 0
transferred to critical care unit | 0
intravenous meropenem | 0
intravenous teicoplanin | 0
severe metabolic acidosis | 0
lactic acidemia | 0
anuria | 0
severe leukopenia | 0
deranged liver function | 0
deranged renal function | 0
deranged coagulation profile | 0
ventricular tachycardia | 12
cardioverted | 12
bradycardia | 12
cardiopulmonary resuscitation | 12
died | 24
blood culture taken | 0
Gram-negative organism | 12
Burkholderia pseudomallei | 12
antibiotic susceptibility testing | 12
polymyxin B minimum inhibitory concentration | 12
antibiogram | 12
VITEK 2 automated system | 12
B. pseudomallei confirmed | 12