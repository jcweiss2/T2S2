76 years old | 0
male | 0
admitted to the hospital | 0
septic arthritis | 0
acute chest pain | 0
chest pain persisted at rest | 0
ECG showed third-degree atrioventricular block | 0
T-waves inversion in inferior leads | 0
lateral ST depressions | 0
triple coronary artery bypass graft (CABG) | -8760
post-myocardial infarction | -8760
left internal mammary artery to left anterior descending artery arterial graft | -8760
saphenous vein grafts (SVGs) aorta (Ao)-circumflex artery | -8760
saphenous vein grafts (SVGs) aorta (Ao)-right coronary artery (RCA) | -8760
coronary angiogram | 1
three patent grafts | 1
aneurysm at the level of the SVG-RCA anastomosis | 1
extravasation of the contrast agent | 1
transthoracic echocardiography | 1
significant pericardial effusion | 1
pericardial effusion compressing the right ventricle | 1
associated haematoma (dry tamponade) | 1
external pacemaker implanted | 1
no invasive mechanical support | 1
pericardiocentesis not performed | 1
admitted to the intensive care unit | 1
transfer to a cardiac surgery centre | 2
passed away from worsening cardiogenic shock | 24
cardiogenic shock | 24 
saphenous vein graft aneurysm post-CABG | -8760 
focal dilatation of the proximal vessel diameter reference | -8760 
aneurysm at the level of the RCA graft | -8760 
asymptomatic | -8760 
choice of percutaneous closure | 1 
surgical management of the aneurysm | 1 
mechanical complications | 1 
fistula | 1 
rupture | 1 
compression of adjacent cardiac or vascular structures | 1 
graft remains patent | 1 
suitable anatomy for stenting | 1 
treated with a covered stent | 1 
balloon occlusion | 1 
coil occlusion | 1 
device occlusion | 1 
loss of RCA perfusion | 1