59 years old | 0
female | 0
lung cancer | -720
pulmonary hypertension | -720
cirrhosis of the liver | -720
hepatitis C positivity | -720
alcohol abuse | -720
consumed raw oysters | -24
generalized lower abdominal pain | -24
admitted to the Emergency Department | 0
non-radiating dull abdominal ache | 0
denied fever | 0
denied chills | 0
no nausea | 0
no vomiting | 0
blood pressure 75/50 mm Hg | 0
pulse rate 100 beats/min | 0
respiratory rate 22 breaths/min | 0
afebrile | 0
temperature 36.7°C | 0
no signs of distress | 0
nontoxic | 0
lungs clear | 0
lower abdominal tenderness | 0
no peritoneal signs | 0
WBC count 0.7 K/uL | 0
hemoglobin level 12.5 g/dL | 0
platelet count 32 K/uL | 0
sodium 144 mEq/L | 0
potassium 3.6 mEq/L | 0
creatinine 1.75 mg/dL | 0
BUN 16 mg/dL | 0
glucose 71 mg/dL | 0
albumin 1.9 g/L | 0
urinalysis positive for infection | 0
+1 protein | 0
+1 blood | 0
+4 urobilinogen | 0
2.5 hyaline casts per high power field | 0
51 to 100 WBCs with clumps | 0
CT scan of the abdomen and pelvis | 0
wall thickening throughout the right colon | 0
inflammation extending along the colon | 0
inflammation surrounding the terminal ileum and appendix | 0
portal venous congestion | 0
pulmonary right lower lobe infiltrate | 0
diagnosis of sepsis with shock | 0
diagnosis of colitis | 0
diagnosis of right lower lobe pneumonia | 0
diagnosis of urinary tract infection | 0
i.v. fluid boluses | 0
norepinephrine | 0
broad-spectrum antibiotics | 0
cefepime | 0
metronidazole | 0
levofloxacin | 0
Granix (tbo-filgrastim) | 0
albuterol/ipratropium nebulization | 0
oxygen saturation above 93% | 0
acute hypoxic respiratory failure | 24
progressive encephalopathy | 24
endotracheal intubation | 24
mechanical ventilation | 24
orogastric tube placement | 24
septic shock | 24
hypotension | 24
albumin administration | 24
sodium bicarbonate infusion | 24
vitamin C sepsis protocol | 24
vitamin C 500 mg i.v. every 8 h | 24
hydrocortisone 100 mg i.v. every 6 h | 24
thiamine 200 mg i.v. every 8 h | 24
doxycycline | 24
blisters and boils on the upper and lower extremities | 30
death | 34
E. tarda in postmortem blood cultures | 34
lung cancer diagnosis | -720
radiation 2 months prior | -720
no chemotherapy | 0
cirrhosis of the liver | -720
iron overload | -720
hemochromatosis | -720
NASH | -720
HCV | -720
obesity | -720