37 years old | 0
    male | 0
    admitted to emergency services | 0
    falling from third floor | 0
    hemodynamically unstable | 0
    aggressive fluid therapy | 0
    X-rays of pelvis | 0
    X-rays of thorax | 0
    chest tube insertion | 0
    pleural effusion | 0
    serosanguineous fluid discharge | 0
    Echo-FAST performed | 0
    abundant free fluid observed | 0
    transferred to operating room | 0
    emergency laparotomy | 0
    hemoperitoneum (4 liters) | 0
    active arterial bleeding | 0
    complete avulsion of hepatic artery | 0
    multiple hepatic lacerations | 0
    remained unstable during surgery | 0
    massive transfusion required | 0
    vasoactive agents required | 0
    ligation of proper hepatic artery | 0
    temporary abdominal closure (vacuum pack) | 0
    admitted to Resuscitation Unit | 0
    hemodynamic recovery | 0
    CT scan performed | 0
    no neurological lesions | 0
    absence of blood flow in hepatic artery | 0
    hepatic dysfunction (ALT 3800) | 0
    hepatic dysfunction (TBil 6) | 0
    hepatic dysfunction (74,000 platelets/μl) | 0
    hepatic dysfunction (IP 40%) | 0
    ischemic hepatitis | 0
    immediate postoperative period | 0
    abdomen closure (definitive) | 72
    bile drainage observed | 168
    suspicion of ischemic cholangiopathy | 168
    poor clinical situation | 168
    transparietohepatic cholangiography performed | 168
    destructuring of bile ducts | 168
    internal-external transhepatic drainage inserted | 168
    clinical improvement | 168
    MRI performed | 168
    multiple hepatic infarctions | 168
    diffuse ischemic cholangiopathy | 168
    septic shock (POD 40) | 960
    cholangitis | 960
    multiple bilomas observed | 960
    irreversible ischemic cholangiopathy | 960
    sepsis control | 960
    multidisciplinary committee decision | 960
    listed for liver transplantation | 960
    liver transplantation performed | 1680
    biliary reconstruction (hepaticojejunostomy) | 1680
    three re-operations post-transplant | 1680
    two arteriographies post-transplant | 1680
    hemoperitoneum post-transplant | 1680
    bilateral mydriasis | 1680
    decreased level of consciousness | 1680
    brain CT scan | 1680
    multiple bilateral ischemic lesions | 1680
    right occipital hemorrhage | 1680
    neurosurgery consultation | 1680
    multidisciplinary session decision | 1680
    therapeutic effort limitation | 1680
    death | 2016
    