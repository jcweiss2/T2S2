73 years old | 0
    male | 0
    prostatectomy | -43800
    prostatic adenocarcinoma | -43800
    Gleason score of 8 (4 + 4) | -43800
    initial protein specific antigen of 17 ng/ml | -43800
    adjuvant radiotherapy | -35064
    hormone therapy | -35064
    acute urine retention | -72
    abdominal pain | -72
    hematuria | -144
    dysuria | -144
    transit disorders | -144
    matter arrest | -144
    decline of general state | -144
    anorexia | -144
    asthenia | -144
    conscious | 0
    asthenic | 0
    performance status at 2 | 0
    diffuse abdominal sensitivity | 0
    painful bladder globe | 0
    bladder catheterization | 0
    venous line administration | 0
    biological check-up | 0
    creatinine at 149 | 0
    K at 6.9 | 0
    blood cells at 14 000/mm3 | 0
    C reactiv protein (CRP) at 450 | 0
    CT scan | 0
    full bladder | 0
    multiple dense formations | 0
    air bubbles | 0
    dense heterogeneous formation at dome | 0
    pneumoperitoneum | 0
    subperitoneal effusion | 0
    hydroaerobic levels | 0
    diffuse mesenteric fat infiltration | 0
    intraperitoneal exploration | 0
    discreet bowel dilatation | 0
    minimal effusion | 0
    hematoma | 0
    bladder breach of ⁓5 cm | 0
    necrotic edges | 0
    inflamed bladder wall | 0
    cystorraphy | 0
    epiploplasty | 0
    Redon drain placement | 0
    renal purification session | 0
    favorable evolution from D1 | 24
    urine clearing | 24
    diuresis of 2400 cc | 24
    Redon to 30 cc | 24
    creatinine at 83 | 24
    K at 5.1 | 24
    blood cells at 11 700/mm3 | 24
    CRP at 324 | 24
    extubated | 48
    recovery of consciousness | 48
    apyretic | 48
    diuresis at 2 L | 48
    Redon removal | 48
    disorder of consciousness | 48
    respiratory distress | 48
    ventricular tachycardia | 48
    cardiorespiratory arrest | 48
    death | 48