57 years old | 0
male | 0
admitted to the hospital | 0
postauricular tingling | -72
discharge-like pain | -72
intense pain | -72
no nausea | -72
no vomiting | -72
no cough | -72
no diarrhea | -72
no limb weakness | -72
no fever | -72
normal physical examination | 0
acupuncture-induced hypersensitivity | 0
normal nervous system examination | 0
normal laboratory examinations | 0
normal coagulation tests | 0
normal thyroid function tests | 0
normal liver and kidney function tests | 0
normal ASO | 0
normal urine analysis | 0
normal stool analysis | 0
normal glycosylated hemoglobin | 0
normal serum homocysteine levels | 0
hypersensitive right lesser occipital nerve | 0
fever | 12
cough | 12
temperature 39.2 °C | 12
pulmonary CT | 24
inflammation in the right lower lung | 24
fine moist rales in the right lower lung | 24
normal oxygen saturation | 24
high fever | 24
respiratory failure | 24
multiple organ failure | 24
bilateral lung infection | 48
wheezing | 48
dyspnea | 48
oxygenation decreased | 48
cyanosis | 48
spots on the trunk and lower extremities | 48
lysin aspirin | 48
noninvasive ventilator-assisted ventilation | 48
imipenem combined with moxifloxacin | 48
oseltamivir | 48
tracheal intubation | 60
hemorrhagic secretions | 60
invasive ventilator | 60
reduced left ventricular systolic and diastolic functions | 60
tolasemide | 60
morphine | 60
metabolic acidosis | 60
sodium bicarbonate | 60
concentrated salt supplementation | 60
noradrenaline | 60
vasoactive dopamine | 60
propofol | 60
midazolam | 60
transferred to ICU | 72
ventilator-assisted ventilation | 72
oxygen saturation 80% | 72
multiple moist rales | 72
heart rate 130 beats/min | 72
strong heart sounds | 72
abdominal softness | 72
borborygmus | 72
vancomycin+biapenem+azithromycin+tami | 72
ECMO treatment | 96
blood oxygen saturation 95% | 96
transfused with red blood cell type A | 96
transfused with plasma | 96
transferred to RICU | 96
nucleic acid PCR for influenza H7N9 virus positive | 96
H7N9 avian influenza virus pneumonia | 96
condition stabilized | 1440
recovered | 2880
discharged | 2880