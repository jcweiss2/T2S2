4.5 years old | 0
male | 0
admitted to the hospital | 0
unconscious | 0
disseminated varicella infection | 0
sepsis | 0
secondary staphylococci infection | 0
transferred to intensive care unit | 0
loss of consciousness | 0
weak spontaneous respiration | 0
intubated | 0
mechanical ventilatory support | 0
death | 96
mild chicken pox | -240
siblings infection | -240
treated with antipyretics | -240
treated with antipruritic lotions | -240
no acyclovir treatment | -240
no vesicular eruption | -240
swelling (right forearm) | -72
bluish discoloration (right forearm) | -72
ulceration (right forearm) | -48
high-grade fever | 0
hypotension | 0
severe dehydration | 0
clear lungs bilaterally | 0
hepatomegaly | 0
abnormal bilateral extensor plantar response | 0
no neck stiffness | 0
excoriated papules (face, trunk, extremities) | 0
serohemorrhagic crusts (face, trunk, extremities) | 0
hemorrhagic necrotic crust (right forearm) | 0
deep ulceration (right forearm) | 0
unremarkable past medical history | 0
high d-Dimer (30 ng/ml) | 0
elevated fibrinogen (465 mg/dl) | 0
prolonged activated partial thromboplastin time (41.6 seconds) | 0
prolonged protrombine time (55 seconds) | 0
elevated white blood cells (9200/mm3) | 0
elevated white blood cells (17,000/mm3) | 24
thrombocytopenia (133,000/mm3) | 0
thrombocytopenia (94,000/mm3) | 24
elevated alanine aminotransferase (324 U/l) | 0
elevated alanine aminotransferase (479 U/l) | 24
elevated aspartate aminotransferase (1402 U/l) | 0
elevated aspartate aminotransferase (1082 U/l) | 24
elevated creatine kinase (35,981 U/l) | 24
elevated CK-MB (1227 U/l) | 24
elevated lactate dehydrogenase (5372 U/l) | 24
elevated sedimantation (42 mm/h) | 24
elevated C-reactive protein (238 mg/l) | 24
urinalysis erythrocytes (5) | 24
urinalysis leukocytes (7) | 24
proteinuria (200 mg/dl) | 24
VZV IgM positive | 0
negative TORCH panel | 0
negative hepatitis markers (HbsAg, anti-HCV) | 0
negative anti-HIV | 0
purpura fulminans | 0
hepatitis | 0
probable rhabdomyolysis | 0
monitorized | 0
vancomycin treatment | 0
cefotaxime treatment | 0
acyclovir treatment | 0
topical silver sulfadiazine cream | 0
hemorrhagic necrotic ulcerative plaque (no expansion) | 96
hemorrhagic necrotic ulcerative plaque (no spread) | 96
