35 years old | 0
woman | 0
diabetes | 0
presented to the emergency department | 0
altered mental status | 0
persistent generalized headache | -168
acetaminophen | -168
ibuprofen | -168
non-productive cough | -96
sore throat | -96
lethargic | -24
confused | -24
unresponsive | -24
random rhythmic movements | -24
no tongue biting | 0
no fecal incontinence | 0
no urinary incontinence | 0
taking food to COVID-19 positive family member | -336
no close contact | -336
no substance use | 0
no smoking | 0
no recent travel | 0
Glasgow Coma Scale 9 | 0
afebrile | 0
temperature 36.6°C | 0
heart rate 93 | 0
blood pressure 133/70 | 0
no nuchal rigidity | 0
negative Brudzinski sign | 0
negative Kernig’s sign | 0
agitation | 0
vomiting | 0
endotracheal intubation | 0
white blood cell count 6900/μL | 0
lactate 1.1 mmol/L | 0
head CT without contrast | 0
no abnormalities on head CT | 0
urinalysis | 0
negative urinalysis | 0
chest x-ray | 0
bilateral patchy infiltrates | 0
nasopharyngeal SARS-CoV-2 PCR positive | 0
pharyngeal swab rapid Streptococcus test positive | 0
Streptococcus pyogenes | 0
blood cultures | 0
vancomycin | 0
ceftriaxone | 0
acyclovir | 0
unsuccessful lumbar puncture | 0
admitted to intensive care unit | 0
fluoroscopy-guided lumbar puncture | 24
cerebrospinal fluid clear then bloody | 24
CSF glucose 109 mg/dL | 24
CSF protein 250 mg/dL | 24
CSF RBC 231/mm3 | 24
CSF WBC 42/mm3 | 24
CSF lymphocytes 62% | 24
CSF monocytes 4% | 24
aseptic meningitis | 24
opening pressure not measured | 24
CSF varicella zoster virus PCR negative | 24
CSF herpes simplex virus 1 PCR negative | 24
CSF herpes simplex virus 2 PCR negative | 24
CSF enterovirus/echovirus PCR negative | 24
CSF syphilis VDRL negative | 24
CSF cryptococcal antigen negative | 24
CSF SARS-CoV-2 testing not performed | 24
MRI brain not performed | 0
C-reactive protein 23.0 mg/L | 0
erythrocyte sedimentation rate 34 mm/hr | 0
D-dimer 0.51 μg/mL | 0
ferritin 125.3 ng/mL | 0
lactate dehydrogenase 267 U/L | 0
interleukin-6 <5 pg/mL | 0
blood cultures negative | 120
CSF cultures negative | 120
vancomycin discontinued | 48
ceftriaxone continued | 0
acyclovir continued | 0
mental status improved | 96
extubated | 96
discharged home | 216
PO penicillin V | 216
PO valacyclovir | 216
