20 years old | 0
female | 0
G1P1 | 0
lactational breast abscess | 0
breastfeeding | -33
pain | -240
erythema | -240
edema | -240
fever | -240
highest temperature 38.3 °C | -240
white blood cell count 14.57 × 10^9/L | -240
neutrophil proportion 83.8% | -240
C-reactive protein 13.76 mg/L | -240
ultrasound showed heterogeneous hypo-echo | -240
antibiotics Amoxicillin Potassium Clavulanate and Metronidazole | -240
symptoms remained poorly controlled | -168
terminate breastfeeding | -168
transferred to hospital | 0
vital signs stable | 0
temperature 36.4 °C | 0
heart rate 105 beats/min | 0
respiratory rate 20 breaths/min | 0
blood pressure 105/69 mmHg | 0
physical exam revealed 8 cm × 6 cm painful mass | 0
ultrasonography showed anechoic mass with internal heterogeneous hypo-echo | 0
white blood cell count 15.43 × 10^9/L | 0
neutrophil proportion 85.3% | 0
CRP 11 mg/L | 0
liver function test normal | 0
renal function test normal | 0
coagulation function test normal | 0
ultrasound-guided needle aspiration failed | 0
milk and pus sent to lab for bacteria test | 0
Cefmetazole administered | 0
body temperature rose to 38.6 °C | 12
surgically removed 150 mL of pus and necrotic tissue | 12
placed 16G indwelling needle for irrigation | 12
placed catheter for drainage | 12
body temperature rose to 41.2 °C | 24
white blood cell count 23 × 10^9/L | 24
neutrophil proportion 96.6% | 24
CRP 138 mg/L | 24
antibiotic changed to Levofloxacin | 24
vital signs deteriorated | 24
heart beat accelerated to 150/min | 24
blood pressure declined to 75/40 mmHg | 24
septic shock | 24
initiated on norepinephrine | 24
transferred to ICU | 24
white blood cell count 40.56 × 10^9/L | 24
neutrophil proportion 97.4% | 24
CRP 186 mg/L | 24
PCT 4.99 | 24
lactic acid 3.98 mmol/L | 24
alkaline phosphatase 164.5 U/L | 24
aspartate aminotransferase 38.7 U/L | 24
alanine aminotransferase 46.3 U/L | 24
albumin 23.7 g/L | 24
total bilirubin 24.1 μmol/L | 24
activated partial thromboplastin time 55.8 s | 24
prothrombin time 24.3 s | 24
INR 2.08 | 24
cultures of blood, stool, and urine samples negative | 24
chest X-ray negative | 24
COVID-19 negative | 24
arterial blood gas analysis showed pH 7.421 | 24
lactic acid 3.98 mmol/L | 24
received treatments including intensive care | 24
placement of central venous catheter | 24
fluid resuscitation | 24
norepinephrine to maintain blood pressure | 24
transfusion of plasma to improve coagulation function | 24
continuous irrigation and drainage of breast abscess | 24
local erythema and edema improved | 48
culture of milk and pus showed Staphylococcal aureus and MRSA | 48
vancomycin prescribed | 48
vitals stable | 120
transferred to department | 120
irrigation and drainage continued | 120
syndrome of erythema, edema and pain disappeared | 168
pus disappeared | 168
drainage extubated | 168
fluid specimen sent to lab for culture | 168
culture revealed no bacteria | 168
discharged | 240
completely asymptomatic during follow-up | 336
completely asymptomatic during follow-up | 480
completely asymptomatic during follow-up | 744