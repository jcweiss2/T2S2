32 years old | 0
white male | 0
started on EPOCH-R | -72
etoposide | -72
vincristine | -72
adriamycin | -72
cyclophosphamide | -72
rituximab | -72
oral prednisone | -72
received Neulasta | -72
rituximab infused | -72
vincristine infused | -72
etoposide infused | -72
adriamycin infused | -72
cyclophosphamide administered | -72
Neulasta administered | -72
first cycle tolerated well | -168
dyspnea | -72
dyspnea worsened with activity | -72
CLS suspected | -72
third cycle without Neulasta | -24
admitted with sudden-onset dyspnea | 0
tachypneic | 0
tachycardic | 0
CT scan negative for pulmonary embolism | 0
diffuse interstitial infiltrate noted | 0
echocardiogram revealed preserved systolic function | 0
no pericardial effusion | 0
started on fluid bolus | 0
administered meropenem | 0
administered vancomycin | 0
worsening respiratory status | 12
transferred to ICU | 12
intubated | 12
started on pressor support | 12
recovered very well | 24
extubated | 48
weaned off pressor support | 48
moved out of ICU | 48
follow-up CT scan revealed bilateral pleural effusion | 72
follow-up CT scan revealed consolidation | 72
continued broad-spectrum antibiotic therapy | 72
possible ventilator-associated pneumonia | 72
Staphylococcus epidermidis growth | 72
positron emission tomography/CT scan confirmed remission of lymphoma | 168
resolution of all abnormalities | 168
completed therapy with CHOP | 168
another 3 cycles | 168
no adverse event | 168
leukocytosis | 0
thrombocytosis | 0
elevated hematocrit | 0
normal BUN | 0
normal creatinine | 0
normal electrolytes | 0
normal liver enzymes | 0
low serum albumin | 0
serum albumin worsened | 48
elevated lactic acid | 0
elevated procalcitonin | 0
exudative pleural effusion | 0
leukocyte count elevated | 0
CLS episode | 0
SCLS | 0
CRS | 0
endothelial dysfunction | 0
noncardiogenic pulmonary edema | 0
hypotension | 0
hypovolemic shock | 0
multi-organ failure | 0
cytokine release | 0
IL-6 trans signaling | 0
endothelial damage | 0
anti-IL-6 strategies | 0
CLS underdiagnosed | 0
avoidance of rituximab therapy | 0
ethical approval not required | 0
informed consent obtained | 0
ORCID iD | 0
