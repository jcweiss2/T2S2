60 years old | 0
male | 0
glomerulonephritis | -672
elevated creatinine | -672
anti-neutrophil cytoplasmic antibody-positive microscopic polyangiitis | -672
methylprednisolone | -72
cyclophosphamide | -72
discharged | -72
nausea | -336
vomiting | -336
diarrhea | -336
intolerance of oral intake | -336
admitted to regional hospital | -336
large volume watery diarrhea | -336
hypovolemic acute kidney injury | -336
hemofiltration | -336
cyclophosphamide reduced | -336
cyclophosphamide ceased | -336
empiric antimicrobial therapy | -336
tazobactam | -336
piperacillin | -336
metronidazole | -336
ganciclovir | -336
secretory diarrhoea | -336
no infective agents identified | -336
vasoactive intestinal polypeptide | -336
chromogranin | -336
diffuse mural thickening of the small and large bowel | -336
denuded and erythematous mucosa | -336
full thickness mucosal ulceration | -336
inflammation | -336
no features of inflammatory bowel disease | -336
no vasculitis | -336
no viral inclusions | -336
diarrhea persisted | 0
antidiarrheals | 0
octreotide | 0
cholestyramine | 0
repeat imaging | 0
repeat stool specimens | 0
repeat endoscopic evaluation | 0
repeat histopathology | 0
regenerative mucosal changes | 0
septic complications | 168
Enterobacter | 168
Candida glabrata | 168
bacteremia | 168
severe acute respiratory distress syndrome | 168
died | 168
post-mortem examination | 168
hemorrhagic ulceration | 168
minimal residual mucosa | 168
no evidence of vasculitis | 168
no evidence of thromboemboli | 168
no definite infectious etiology | 168
herpes simplex virus-1 DNA | 168
diffuse alveolar damage | 168
metastatic pulmonary calcification | 168
Enterobacter faecium | 168
Candida krusei | 168
Pneumocystis jiroveci | 168
inflammatory bowel disease | -672
neutropenic typhilitis | -336
auto-immune | -336
vasculitic | -336
infective colitis | -336
carcinoid syndrome | -336
ischemic bowel | -336
prophylactic antibiotics | 0
prophylactic antivirals | 0
prophylactic antifungals | 0
intravenous fluids | 0
electrolytes | 0
total parenteral nutrition | 0
glucocorticoids | 0
infliximab | 0
intestinal transplantation | 168