54 years old | 0
female | 0
height 170 cm | 0
weight 68 kg | 0
heavy smoker | 0
no drug allergy | 0
bilateral cataract extraction | -8760
breast augmentation | -8760
abdominoplasty | -8760
admitted to hospital | 0
screening gastroscopy | 0
colonoscopy | 0
sedation | 0
oxygen supplementation | 0
meperidine | 0
midazolam | 0
propofol | 0
gastroscopy started | 0
bradycardia | 10
asystole | 10
premature ventricular contraction | 10
bizarre QRS wave | 10
undetectable blood pressure | 10
xylocaine | 10
atropine | 10
epinephrine | 10
hydrocortisone | 10
face mask ventilation | 10
sinus tachycardia | 10
systemic blood pressure improved | 10
regained consciousness | 10
acute chest pain | 10
pulmonary edema | 10
dyspnea | 10
hypoxia | 10
procedure aborted | 10
transferred to ICU | 10
EKG | 10
chest X-ray | 10
diffuse bilateral infiltrations | 10
transthoracic echocardiography | 10
global hypokinesia | 10
ejection fraction 20-29% | 10
respiratory acidosis | 10
ABGs | 10
Lasix | 10
dobutamine | 10
improved clinically | 12
saturation improved | 12
BiPAP | 12
weaning of dobutamine started | 24
troponin level 0.08 | 0
troponin level 0.54 | 12
troponin level 0.58 | 18
coronary angiography | 24
no significant coronary stenosis | 24
fully recovered | 48
discharged | 96
carvedilol | 96
rabeprazole sodium | 96
follow-up | 2160