48 years old | 0
non-alcoholic | 0
non-smoker | 0
female | 0
presented to out-hospital clinic | -168
cough | -168
generalized myalgia | -168
arthralgia | -168
fever | -168
physical examination | 0
temperature 36.9°C | 0
pulse 76/m | 0
blood pressure 132/78 mmHg | 0
oxygen saturation 96% | 0
body mass index 26 | 0
diffuse arthralgia | 0
myalgia | 0
no previous medical history | 0
no chronic diseases | 0
no previous treatment | 0
no family history | 0
elevated erythrocyte sedimentation rate | 0
elevated C-reactive protein | 0
elevated creatine kinase | 0
nasopharyngeal swab confirmed COVID-19 | 0
mild disease (WHO classification) | 0
computed tomography pulmonary infiltrations | 0
hospitalized in COVID-19 isolation | 0
admitted to ICU | 72
confusion | 72
high fever 39.8°C | 72
tachycardia 125/m | 72
hypotension 75/40 mmHg | 72
Glasgow score 10/15 | 72
white blood cells 10,000 | 72
erythrocyte sedimentation rate 61 m/h | 72
C-reactive protein 36 mg/dl | 72
creatine phosphokinase 542310 IU | 72
myoglobin >15,000 g/l | 72
aspartate aminotransferase 1246 U/L | 72
alanine aminotransferase 986 U/L | 72
urea 154 | 72
creatinine 2.8 | 72
normal troponin | 72
normal D-dimer | 72
treated with oxygen 12 l/min | 72
intravenous normal saline | 72
bicarbonate 1.4% | 72
epinephrine | 72
azithromycin | 72
methyl prednisone 250 mg IV | 72
enoxaparine 4000 IU SC | 72
intubated | 72
mechanically ventilated | 72
dialysis therapy | 72
anuria | 72
metabolic acidosis | 72
hyperkalemia | 72
died | 96
cardiac arrest | 96
hemodynamic deterioration | 96
rhabdomyolysis | 0
musculoskeletal manifestations (fatigue, myalgia, arthralgia, etc.) | 0
dark red or brown urine | 0
decreased urination | 0
abdominal pain | 0
muscle pain | 0
lack of consciousness | 0
acute renal failure | 72
disseminated intravenous coagulation | 72
48 years old| 0
non-alcoholic| 0
non-smoker| 0
female| 0
presented to out-hospital clinic| -168
cough| -168
generalized myalgia| -168
arthralgia| -168
fever| -168
physical examination| 0
temperature 36.9°C| 0
pulse 76/m| 0
blood pressure 132/78 mmHg| 0
oxygen saturation 96%| 0
body mass index 26| 0
diffuse arthralgia| 0
myalgia| 0
no previous medical history| 0
no chronic diseases| 0
no previous treatment| 0
no family history| 0
elevated erythrocyte sedimentation rate| 0
elevated C-reactive protein| 0
elevated creatine kinase| 0
nasopharyngeal swab confirmed COVID-19| 0
mild disease (WHO classification)| 0
computed tomography pulmonary infiltrations| 0
hospitalized in COVID-19 isolation| 0
admitted to ICU| 72
confusion| 72
high fever 39.8°C| 72
tachycardia 125/m| 72
hypotension 75/40 mmHg| 72
Glasgow score 10/15| 72
white blood cells 10,000| 72
erythrocyte sedimentation rate 61 m/h| 72
C-reactive protein 36 mg/dl| 72
creatine phosphokinase 542310 IU| 72
myoglobin >15,000 g/l| 72
aspartate aminotransferase 1246 U/L| 72
alanine aminotransferase 986 U/L| 72
urea 154| 72
creatinine 2.8| 72
normal troponin| 72
normal D-dimer| 72
treated with oxygen 12 l/min| 72
intravenous normal saline| 72
bicarbonate 1.4%| 72
epinephrine| 72
azithromycin| 72
methyl prednisone 250 mg IV| 72
enoxaparine 4000 IU SC| 72
intubated| 72
mechanically ventilated| 72
dialysis therapy| 72
anuria| 72
metabolic acidosis| 72
hyperkalemia| 72
died| 96
cardiac arrest| 96
hemodynamic deterioration| 96
rhabdomyolysis| 0
musculoskeletal manifestations (fatigue, myalgia, arthralgia, etc.)| 0
dark red or brown urine| 0
decreased urination| 0
abdominal pain| 0
muscle pain| 0
lack of consciousness| 0
acute renal failure| 72
disseminated intravenous coagulation| 72
