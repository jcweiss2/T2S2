77 years old | 0
female | 0
breast cancer | -6720
chemotherapy | -6720
radiation to the chest | -6720
severe aortic stenosis | -6720
coronary artery disease | -6720
90% occlusion of the left anterior descending artery | -6720
admitted to the hospital | 0
tissue aortic valve replacement | 0
saphenous vein graft bypass | 0
midline sternotomy | 0
induction of anesthesia | 0
intubation | 0
dissection of the left internal mammary artery | 0
atretic left internal mammary artery | 0
use of the greater saphenous vein | 0
small greater saphenous vein | 0
decline in cerebral head saturations | 0
reduced mean arterial perfusion | 0
reduced cerebral artery perfusion | 0
use of vasopressors | 0
extubation | 2
persistent lactic acidosis | 2
high-dose vasopressor support | 2
mixed cardiogenic and vasoplegic shock | 2
lethargy | 15
leftward gaze | 15
right upper extremity weakness | 15
resolution of symptoms | 15
tongue ecchymoses | 15
tongue numbness | 15
dysgeusia | 15
CT scan of the head | 15
no acute hemorrhage | 15
CT angiogram of the brain and neck | 15
no large vessel occlusion | 15
mild calcification at the bifurcation of the right common carotid artery | 15
50% focal stenosis of the distal left common carotid artery | 15
completely occluded right lingual artery | 15
mild distal collateral flow | 15
multifocal irregularities of the left lingual artery | 15
normal postoperative platelet count | 15
normal prothrombin time | 15
normal international normalized ratio | 15
normal fibrinogen | 15
no prior history of known vasculitic disease | 15
normal ADAMTS13 inhibitor screen | 15
volume resuscitation | 15
low-dose epinephrine | 15
high-dose norepinephrine | 15
high-dose vasopressin | 15
improvement of systemic vascular resistance | 48
otolaryngology service consultation | 48
serial examinations of the patient’s tongue | 48
evaluation with multiple flexible bronchoscopes | 48
persistent tongue numbness | 48
persistent dysgeusia | 48
supportive therapy | 48
improvement of symptoms | 48
return of tongue sensation | 1440
return of taste | 1440
discharge from the hospital | 1440