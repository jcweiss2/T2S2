58 years old | 0
male | 0
fever | -168
fatigue | -168
cough | -168
severe shortness of breath | -168
oxygen saturation of 70% | 0
intubated | 0
bilateral diffuse pulmonary infiltrates | 0
interstitial thickening | 0
bilateral basal consolidation | 0
PCR nasopharyngeal swab positive for SARS-CoV-2 | 0
pancytopenia | 0
white blood cell count 2.6 × 103/μL | 0
absolute neutrophil count 1.8 × 103/μL | 0
hemoglobin 12.1 g/dL | 0
platelet count 85 × 103/μL | 0
acute kidney injury | 0
serum creatinine level 120 μmol/L | 0
transaminitis | 0
alanine aminotransferase 170.2 U/L | 0
aspartate aminotransferase 330 U/L | 0
lactic acid dehydrogenase 857 U/L | 0
hydroxychloroquine 400 mg | 0
azithromycin 500 mg | 0
interleukin-6 1,843 pg/mL | 0
D-dimer 73.37 mg/L | 0
ferritin 2,166.0 μg/L | 0
cytokine storm | 0
tocilizumab 400 mg | 0
methylprednisone 40 mg | 0
intravenous immunoglobulin 0.4 g/kg | 0
severe sepsis | 0
vasopressors | 0
broad-spectrum antibiotics | 0
antifungals | 0
sustained low-efficiency dialysis | 0
ultrasound abdomen normal spleen | 0
granulocyte colony-stimulating factor | 0
persistent pancytopenia | 384
white blood cell count 0.5 × 103/μL | 384
absolute neutrophil count 0.3 × 103/μL | 384
hemoglobin 8.4 g/dL | 384
platelet count 74 × 103/μL | 384
peripheral blood smear pancytopenia | 384
red cell agglutination | 384
atypical lymphoid cells | 384
hairy cells | 384
monocytopenia | 384
bone marrow aspirate hypocellular | 384
decreased trilineage hematopoiesis | 384
bone marrow core biopsy hypercellular | 384
infiltration with atypical cells | 384
decreased erythropoiesis | 384
decreased granulopoiesis | 384
increased megakaryocytes | 384
increased histiocytes | 384
hemosiderin-laden macrophages | 384
reticulin fibrosis | 384
CD20 positivity | 384
DBA.44 positivity | 384
PAX5 positivity | 384
annexin A1 positivity | 384
cyclin D1 positivity | 384
CD25 positivity | 384
V600E-mutant BRAF protein positivity | 384
flow cytometry monotypic B cells | 384
CD45 positivity | 384
CD19 positivity | 384
CD79b positivity | 384
FMC7 positivity | 384
CD11c positivity | 384
CD103 positivity | 384
CD10 positivity | 384
CD200 positivity | 384
cBCL2 positivity | 384
IgM positivity | 384
lambda light chain restriction | 384
CD23 negativity | 384
CD5 negativity | 384
CD123 negativity | 384
CD38 negativity | 384
CD43 negativity | 384
IgD negativity | 384
FISH analysis normal | 384
cytogenetic analysis normal male karyotype | 384
BRAF V600 mutation confirmed | 384
diagnosis of hairy cell leukemia | 384
absence of splenomegaly | 0
lack of CD123 expression | 384
expression of CD10 | 384
decision to wait for COVID-19 recovery | 384
