33 years old | 0
diabetic | 0
male | 0
presented to the emergency department | 0
left thigh pain | 6
pain woke him up from sleep | 6
pain not relieved with over-the-counter medication | 6
denied history of recent trauma | 0
former smoker | -336
quit smoking | -336
denied personal history of hypercoagulable disorders | 0
denied family history of hypercoagulable disorders | 0
denied illicit substance use | 0
review of systems was negative | 0
lack of respiratory symptoms | 0
diffusely swollen left thigh | 0
cyanotic left thigh | 0
tender left thigh | 0
tense left thigh | 0
no evidence of trauma | 0
left leg cool to touch | 0
intact motor function | 0
intact sensory function | 0
soft left calf | 0
palpable femoral pulse | 0
popliteal artery signal present | 0
posterior tibial artery signal present | 0
soft right lower extremity compartments | 0
palpable femoral pulse (right) | 0
palpable popliteal pulse (right) | 0
palpable dorsalis pedis pulse (right) | 0
palpable posterior tibial pulse (right) | 0
computed tomography angiography performed | 0
bilateral multifocal ground-glass opacities | 0
consolidation in lower lobes | 0
concerning for COVID-19 infection | 0
acute occlusion of left mid-superficial femoral artery | 0
no evidence of reconstitution | 0
significant left thigh musculature swelling | 0
therapeutic anticoagulation with unfractionated heparin | 0
taken to operating room | 0
angiography of lower extremity | 0
fasciotomy of left thigh | 0
angiogram through right transfemoral approach | 0
no arterial thrombosis | 0
contiguous sluggish flow to foot | 0
elevated anterior compartment pressures | 0
elevated posterior compartment pressures | 0
decompressive fasciotomy of two compartments | 0
lateral thigh incision | 0
healthy left thigh muscles | 0
pink muscles | 0
contractile muscles | 0
venous duplex ultrasound negative for deep venous thrombosis | 0
normal arterial flow on angiography | 0
suspected viral myositis in COVID-19 | 0
kept on full-dose anticoagulation | 0
concern for hypercoagulable state | 0
unremarkable muscle biopsy | 0
admitted to intensive care unit | 0
fully anticoagulated | 0
empirical COVID-19 treatment with hydroxychloroquine | 0
empirical COVID-19 treatment with azithromycin | 0
awaiting PCR results | 0
positive PCR test | 0
negative hypercoagulable workup | 0
normal creatine kinase on admission | 0
creatine kinase remained normal until postoperative day 9 | 216
improved after initial operation | 0
improved left thigh | 0
nonedematous left calf | 0
no respiratory symptoms during hospitalization | 0
acute left calf pain on postoperative day 9 | 216
elevated compartment pressures | 216
palpable distal pulses | 216
no concern for arterial thrombosis | 216
emergent four-compartment fasciotomy | 216
significantly edematous muscle | 216
deteriorated clinical condition | 216
developed diabetic ketoacidosis | 216
developed acute kidney injury | 216
developed thrombocytopenia | 216
platelet count 19,000/μL | 216
developed bilateral subsegmental pulmonary embolism | 216
developed bilateral iliofemoral thrombosis | 216
developed inferior vena cava thrombosis | 216
developed diffuse arterial thrombosis (right femoropopliteal) | 216
developed diffuse arterial thrombosis (left infrapopliteal) | 216
cold extremities bilaterally | 216
intact motor function | 216
intact sensory function | 216
unsafe to attempt surgery | 216
maintained on anticoagulation | 216
right calf pain on postoperative day 11 | 264
elevated compartment pressures | 264
improved clinical course | 264
demarcation at toes bilaterally | 264
revascularization not attempted | 264
taken to operating room | 264
right lower extremity four-compartment fasciotomy | 264
edematous muscle | 264
dusky muscle | 264
right thigh compartment syndrome on postoperative day 13 | 312
taken to operating room | 312
three-compartment fasciotomy | 312
compartment syndrome due to arterial and venous thrombosis | 312
remained on therapeutic anticoagulation | 312
prophylactic broad-spectrum antibiotics | 312
received convalescent antibody plasma therapy on postoperative day 16 | 384
left below-knee amputation | 384
right above-knee amputation | 384
demarcation of lower extremities | 384
discharged to rehabilitation facility | 384
elevated D-dimer | 0
elevated C-reactive protein | 0
proinflammatory state | 0
hypercoagulable state | 0
