50 years old | 0
male | 0
admitted to the hospital | 0
unsteady gait | -72
weakness | -72
somnolence | -72
systolic heart failure | -6720
ejection fraction of 21% | -6720
remote orthotopic liver transplantation | -6720
alcohol- and hepatitis C-induced cirrhosis | -6720
acute renal failure | -6720
hemodialysis | -6720
nonadherence to immunosuppressant medications | -336
tacrolimus | -336
everolimus | -336
creatinine of 6.1 mg/dL | 0
blood urea nitrogen of 23 mg/dL | 0
prothrombin time of 15.9 seconds | 0
partial thromboplastin time of 35 seconds | 0
international normalized ratio of 1.5 | 0
leukocytosis of 13.4 × 10^9/L | 0
paracentesis | 0
bloody ascitic fluid | 0
no evidence of spontaneous bacterial peritonitis | 0
vancomycin | 0
piperacillin/tazobactam | 0
hypotensive to 73/35 mm Hg | 12
hemoglobin dropped from 7.4 to 5.6 gm/dL | 12
packed red blood cells | 12
Ringer's lactate | 12
albumin | 12
fresh frozen plasma | 12
hemoglobin improved to 7.1 mg/dL | 12
hemodynamics normalized | 12
computed tomography of the abdomen and pelvis | 12
intraperitoneal active extravasation | 12
injury to the right inferior epigastric artery or an intercostal artery | 12
interventional radiology fluoroscopy suite | 24
right common femoral artery accessed | 24
wire advanced centrally | 24
5Fr sheath placed | 24
Mikaelson catheter | 24
right 10th, 11th, and 12th intercostal arteries selected | 24
arteriograms | 24
embolization of the right 11th and 12th intercostal arteries | 24
gelatin foam | 24
completion angiogram | 24
hemoglobin decreased to 5.6 mg/dL | 48
repeat computed tomography of the abdomen and pelvis | 48
persistent arterial extravasation | 48
additional packed red blood cells | 48
platelets | 48
fresh frozen plasma | 48
prothrombin complex concentrate | 48
conservative management | 48
critical care team discussion | 48
interventional radiology team discussion | 48
surgical team discussion | 48
Doppler ultrasound | 72
color jet extending into the distended peritoneum | 72
thrombin injection | 72
bovine thrombin | 72
thrombin-saline mixture | 72
vascular jet no longer visualized | 72
hemoglobin remained stable | 72
hemodynamics improved | 72
persistent leukocytosis | 96
systemic inflammatory response syndrome | 96
no identified source of infection | 96
empiric vancomycin and piperacillin/tazobactam | 96
immunosuppressant medications restarted | 96
transferred to outside hospital | 120