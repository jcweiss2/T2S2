63 years old | 0
female | 0
alcohol use disorder | 0
type 2 diabetes mellitus | 0
hypertension | 0
chronic pancreatitis | 0
pseudocyst | 0
admitted to the ICU | 0
mixed hemorrhagic/distributive shock | 0
acute gastrointestinal bleed | 0
diabetic ketoacidosis | 0
lethargic | -24
declining responsiveness | -24
hypothermic | -24
hypotensive | -24
hemoglobin of 13 g/dL | -24
glucose greater than 1500 mg/dL | -24
beta-hydroxybutyrate greater than 22.50 mmol/L | -24
creatinine of 3.55 mg/dL | -24
blood urea nitrogen (BUN) of 101 mg/dL | -24
bicarbonate of 5 mmol/L | -24
pH of 7.01 | -24
hematemesis | -24
intubation | -24
placement of a right internal jugular vein central line | -24
insulin drip | -24
pantoprazole drip | -24
ceftriaxone | -24
transfer to hospital | -24
afebrile | 0
tachycardic | 0
norepinephrine infusion | 0
vasopressin infusion | 0
pH of 7.21 | 0
bicarbonate of 22 mmol/L | 0
glucose of 902 mg/dL | 0
anion gap of 28 mmol/L | 0
potassium of 3.7 mmol/L | 0
BUN of 84 mg/dL | 0
creatinine of 2.47 mg/dL | 0
lipase of 69 U/L | 0
C-reactive protein of 262 mg/L | 0
sedimentation rate of greater than 120 mm/h | 0
undetectable ethanol | 0
hemoglobin of 15 g/dL | 0
platelets of 165 000 per cu mm | 0
white blood cell count of 3300 per cu mm | 0
infectious diseases workup | 0
blood cultures | 0
sputum cultures | 0
urine cultures | 0
chest X-ray | 0
broad-spectrum antimicrobial coverage | 0
piperacillin/tazobactam | 0
Candida species in blood cultures | 24
micafungin | 24
C. albicans | 24
line holiday | 48
removal of arterial line | 48
removal of right internal jugular vein central line | 48
transthoracic echocardiogram | 48
CT of the chest | 48
CT of the abdomen and pelvis | 48
ophthalmologic exam | 48
plain films of left hip | 48
hip aspiration | 48
upper and lower extremity duplexes | 120
deep vein thrombus (DVT) in the right internal jugular vein | 120
heparin drip | 120
clearance of clot and blood cultures | 144
fluconazole | 144
enoxaparin | 144
discharge to a skilled nursing facility | 744
Candida thrombophlebitis | 120
septic thrombophlebitis | 120
infected thrombi | 120
fungemia | 24
sepsis | 0
organ dysfunction | 0
mechanical ventilation | 0
Candida colonization | 0
broad-spectrum antibiotic exposure | 0
arterial or central venous catheter | 0
new-onset sepsis | 0
empiric coverage with micafungin | 0
invasive fungal infection-free survival | 0