48 years old | 0
male | 0
incarcerated | 0
admitted to the hospital | 0
multisystem sarcoidosis | -672
bone marrow involvement | -672
liver involvement | -672
lymph nodes involvement | -672
non-caseating granulomas | -672
progressive abdominal pain | -2304
100-pound weight loss | -2304
nausea | -2304
vomiting | -2304
paraplegia | -5184
urinary retention | -5184
asthma | 0
type 2 diabetes mellitus | 0
gastroesophageal reflux disease | 0
hiatal hernia | 0
hypertension | 0
alcoholism | 0
magnetic resonance imaging (MRI) of the thoracic spine | -2592
degenerative disc disease of the thoracic spine | -2592
MRI of the lumbar spine | -2592
disc bulging at L5–S1 | -2592
albuterol | -672
terazosin | -672
oxybutynin | -672
pantoprazole | -672
admitted to an outside hospital | -672
diagnosed with sarcoidosis | -672
weight loss | -672
abdominal pain | -672
leukopenia | -672
anemia | -672
computed tomography (CT) abdomen and pelvis | -672
large mesenteric and retroperitoneal lymph node adenopathy | -672
splenomegaly | -672
large splenic masses | -672
heterogenous liver parenchyma | -672
liver biopsy | -672
bone marrow biopsy | -672
retroperitoneal lymph node biopsy | -672
non-necrotizing granulomatous inflammation | -672
necrotizing granulomatous inflammation | -672
prednisone | -672
methotrexate | -672
admitted to the same hospital | -72
chest pain | -72
anorexia | -72
nausea | -72
vomiting | -72
abdominal pain | -72
hypotensive | -72
blood pressure 85/63 mmHg | -72
temperature 98.6°F | -72
pulse 117 beats per minute | -72
respiratory rate 22 breaths per minute | -72
oxygen saturation 95% | -72
CT thorax | -72
moderate right and small-to-moderate left pleural effusions | -72
CT abdomen and pelvis | -72
stable changes | -72
new moderate ascites | -72
urine and blood cultures | -72
lactate 2.3 mmol/L | -72
INR >12 | -72
fibrinogen 50 mg/dL | -72
ALT 86 IU/L | -72
AST 204 IU/L | -72
white blood cell count (WBC) 0.8 K/uL | -72
hemoglobin (Hb) 7.9 g/dL | -72
platelets 92 K/uL | -72
admitted to the Intensive Care Unit (ICU) | -72
suspected sepsis | -72
intravenous fluids | -72
cefepime | -72
vancomycin | -72
Vitamin K | -72
Hematology | -72
Infectious Disease | -72
Rheumatology | -72
cefepime and vancomycin stopped | -48
methylprednisolone | -48
transferred to our hospital | 0
bone marrow biopsy | 24
hypocellular bone marrow | 24
trilineage hematopoiesis | 24
no malignancy | 24
no granulomas | 24
occasional histiocytic hemophagocytosis | 24
soluble CD 25 (soluble interleukin-2 receptor) | 24
elevated at 70 000 pg/mL | 24
etoposide | 48
IVIG | 48
ferritin improved | 72
kidney function worsened | 72
creatinine 1.26 mg/dL to 3.34 mg/dL | 72
second dose of etoposide decreased | 96
vancomycin discontinued | 96
Sustained Low Efficiency Dialysis (SLED) | 120
bumetanide | 120
obtunded | 144
hypotensive | 144
hypothermic | 144
intubated | 144
lactic acidosis | 144
ALT 1985 IU/L | 144
AST 3322 IU/L | 144
LDH 10,692 IU/L | 144
haptoglobin <30 mg/dL | 144
ferritin 65,620 ng/ml | 144
lactate 14 mmol/L | 144
WBC 0.1 K/uL | 144
hemoglobin 6.5 | 144
platelets <10 k/uL | 144
ANC 0 k/uL | 144
GI bleed | 144
hypovolemic and hemorrhagic shock | 144
intracranial hemorrhage | 144
CT head | 144
no evidence of intracranial hemorrhage | 144
pulseless electrical activity arrest | 168
resuscitation efforts unsuccessful | 168
died | 168