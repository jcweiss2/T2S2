52 years old | 0
female | 0
admitted | 0
fever | -240
cough | -240
breathlessness | -240
progressive dyspnea | -240
decrease urine output | -240
no history of abdominal pain | 0
no history of dysuria | 0
no history of trauma | 0
no recent use of non-steroidal anti-inflammatory medication | 0
breathless | 0
blood pressure 150/90 mmHg | 0
temperature 40°C | 0
respiratory rate 30 breaths/min | 0
heart rate 100 bpm | 0
hemoglobin 10.3 g/l | 0
total white cell count 9.88 × 103/μl | 0
neutrophils 74% | 0
lymphocytes 20% | 0
monocytes 4% | 0
eosinophils 2% | 0
platelet count 211 × 103/μl | 0
serum creatinine 10.8 mg/dl | 0
sodium 138 mEq/l | 0
potassium 5.3 mEq/l | 0
blood urea 76 mg/dl | 0
blood glucose 72 mg/dl | 0
renal ultrasound normal sized kidneys | 0
hyper reflective cortex | 0
serological tests negative for malaria | 0
serological tests negative for leptospirosis | 0
serological tests negative for dengue | 0
serological tests negative for viral hepatitis | 0
initial blood cultures sterile | 0
initial urine cultures sterile | 0
initial sputum cultures sterile | 0
urinalysis proteinuria | 0
urinalysis hematuria | 0
two to five fine granular casts | 0
SCr phosphokinase levels unremarkable | 0
liver function test chest radiograph unremarkable | 0
antinuclear antibody negative | 0
anti-double-stranded deoxyribonucleic acid negative | 0
anti-neutrophil cytoplasmic antibody negative | 0
anti-globular basement membrane antibody negative | 0
coombs’ test negative | 0
cryoglobulins negative | 0
C-reactive protein negative | 0
complement components (C3 and C4) low | 0
HIV negative | 0
hepatitis B surface antigen negative | 0
hepatitis C virus negative | 0
influenza H1N1 virus detected | 0
exposure to swine flu positive patient | 0
oseltamivir | 0
antibiotic | 0
fluid replacement | 0
dialysis | 0
peritoneal dialysis | 0
oliguric | 0
required intermittent hemodialysis | 0
hemodialysis 5 times | 0
temporary jugular dialysis catheter | 0
renal biopsy mesangial proliferative glomerulonephritis | 0
acute tubule interstitial nephritis | 0
methyl prednisolone 500 mg | 0
oral prednisolone 1 mg/kg/day | 0
discharged | 0
SCr 1.5 mg/dl | 0
SCr 1 mg/dl at 1 month follow-up | 720
