75 years old | 0  
    male | 0  
    admitted via casualty | 0  
    collapse secondary to seizures | 0  
    intermittent dialysis for end stage renal disease (ESRD) | 0  
    left lacunar infarct in temporal lobe | 0  
    coronary artery bypass graft (CABG) in 2000 | 0  
    hypertension | 0  
    chronic obstructive pulmonary disease (COPD) | 0  
    atrial fibrillation | 0  
    warfarin | 0  
    confused | 0  
    both pupils equal | 0  
    reactive to light | 0  
    Glasgow coma scale of 12/15 | 0  
    tachycardic | 0  
    hypotensive | 0  
    tachypnoeic | 0  
    raised renal parameters | 0  
    altered coagulation profile | 0  
    electrocardiogram | 0  
    computed tomography (CT) of brain | 0  
    no new changes on CT of brain | 0  
    deterioration | 0  
    intubated | 0  
    mechanically ventilated | 0  
    right radial artery cannulated | 0  
    blood pressure monitoring | 0  
    ABG measurements | 0  
    cannulation remained in situ for 7 days | 0  
    cannulation removal | 168  
    inflammation at skin site 5 days post-removal | 168  
    wound swab grew MRSA | 168  
    inflammation appeared to settle | 168  
    distinct bulging of radial artery 8 days later | 312  
    ultrasound performed | 312  
    radial artery pseudoaneurysm diagnosed | 312  
    angiogram confirmation | 312  
    radial artery compression as treatment | 312  
    rupture after a week | 384  
    surgical intervention | 384  
    surgical exploration confirmed 6x5 cm pseudoaneurysm | 384  
    MRSA infection | 168  
    catheter-related sepsis risk factors | 0  
    duration of catheterization (7 days) | 0  
    age (75 years old) | 0  
    ESRD on dialysis | 0  
    anticoagulation with warfarin | 0  
    hypotension | 0  
    multiple attempts (3) during cannulation | 0  
    no external signs of infection at cannulation site | 0  
    hospital protocol for cannula change | 0  
    use of ultrasound for cannulation in high-risk patients | 0  
    aseptic precautions | 0  
    immunocompromised state | 0  
    percutaneous injection of bovine thrombin under ultrasound guidance | 384  
    mechanical compression | 384  
    micro vascular surgeries | 384  