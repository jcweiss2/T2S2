73 years old | 0
male | 0
South Asian ethnicity | 0
progressive chronic kidney disease | 0
obstructive uropathy | 0
recurrent urosepsis | 0
hydronephrotic left kidney | 0
insertion of J-J ureteric stent | -15864
type 2 diabetes mellitus | 0
ischaemic heart disease | 0
myocardial infarction | -16224
hypertension | 0
no history of cardiac dysrhythmia | 0
no prothrombotic diathesis | 0
no cerebrovascular disease | 0
no family history of renal disease | 0
no family history of cerebrovascular disease | 0
not on maintenance antiplatelet agents | 0
not on oral anticoagulants | 0
non-smoker | 0
no alcohol consumption | 0
emergency admission to intensive care unit | -1800
pulmonary oedema | -1800
oliguria | -1800
serum creatinine 10.2 mg/dL | -1800
maintenance thrice weekly HD via right internal jugular tunnelled cuffed central venous catheter | -1800
acute stroke presentation | 0
acute right hemiparesis | 0
aphasia | 0
duration of 90 minutes | 0
routine HD 24 hours prior | -24
blood pressure 190/87 mmHg | 0
capillary blood glucose 86.5 mg/dL | 0
Glasgow Coma Score 15/15 | 0
sinus rhythm on electrocardiogram | 0
urgent CT scan of brain | 0
acute ischaemic stroke affecting superior parasagittal cortex of left frontal lobe | 0
no evidence of intracranial haemorrhage | 0
transferred to local acute stroke centre | 0
blood pressure 176/75 mmHg | 0
mild right facial droop | 0
right hemiparesis | 0
power 3/5 in upper limb | 0
power 0/5 in lower limb | 0
increased muscle tone in upper limb | 0
lower limb hyper-reflexia | 0
upgoing plantar response in lower limb | 0
dysphasia with receptive and expressive elements | 0
no cardiac murmurs | 0
no carotid bruits | 0
clinically euvolaemic | 0
NIH stroke score 8 | 0
no absolute contraindications to thrombolysis | 0
eligible for trial enrolment | 0
informed consent | 0
received 54 mg rtPA | 240
repeat CT brain scan | 264
small area of haemorrhagic transformation within original infarct | 264
no other interval change | 264
clinically stable | 264
required sodium valproate | 264
required clobazam | 264
intermittent left upper limb myoclonus | 264
responded well to therapy | 264
echocardiography revealed borderline left ventricular hypertrophy | 264
24-hour Holter during interdialytic period | 264
sinus rhythm | 264
1-hour paroxysm of asymptomatic atrial fibrillation | 264
terminated spontaneously | 264
no significant carotid stenosis | 264
transferred to specialist renal stroke rehabilitation unit | 96
inpatient for following month | 96
upper limb power improved to 4/5 proximally | 96
upper limb power improved to 3/5 distally | 96
lower limb power improved to 4/5 proximally | 96
dysphasia improved | 96
residual mild expressive deficit | 96
discharged home | 840
remains stable on maintenance HD | 840
