85 years old | 0
male | 0
admitted to the hospital | 0
skin ulceration | 0
left upper limb | 0
lethargy | 0
fever | -24
stabbed in the left upper limb | -24
drowsiness | -24
maximum body temperature of 38.8 °C | -24
skin in the left upper limb was ulcerated | 0
red and swollen | 0
petechiae | 0
ecchymosis | 0
White blood cell count (WBC) 11.77 × 10^9/L | 0
procalcitonin (PCT) > 100 ng/mL | 0
lactate (Lac) 4.28 mmol/L | 0
cultures of blood | 0
secretions | 0
fluid seeping from the broken blisters | 0
antibiotic sensitivity test | 0
metagenomic analysis of pathogens in blood sample | 0
next-generation sequencing (NGS) | 0
anti-infection treatment | 0
azithromycin | 0
tienam | 0
rehydration | 0
pressure promotion | 0
anticoagulation | 0
admitted to the emergency intensive care unit (EICU) | 24
septic shock | 24
diabetes | -7200
alcoholism | -7200
meropenem | 24
levofloxacin | 24
norepinephrine | 24
vasopressin | 24
argatroban | 24
ulinastatin | 24
multiple incisions | 24
decompression | 24
drainage | 24
gentamicin | 24
magnesium sulfate | 24
tracheal intubation | 24
ventilator | 24
fever | 48
ulceration | 48
oedema | 48
improvement | 48
new petechiae | 48
tension blisters | 48
dark purple skin | 48
patchy ecchymosis | 48
doxycycline | 48
blood culture identification | 72
antibiotic sensitivity test | 72
V. vulnificus | 72
liver function reexamination | 96
alanine aminotransferase (ALT) level of 2295 U/L | 96
aspartate aminotransferase (AST) level of 1273 U/L | 96
discontinued doxycycline | 96
body temperature was normal | 192
skin ulceration alleviated | 192
redness alleviated | 192
WBC 9.09 × 10^9/L | 192
PCT 2.68 ng/mL | 192
Lac 1.74 mmol/L | 192
ALT 281 U/L | 192
AST 44 U/L | 192
sedation stopped | 192
spontaneous breathing trial (SBT) | 192
extubated | 192
noninvasive ventilator-assisted ventilation | 192
no fever | 408
vital signs stable | 408
swelling improved | 408
ulceration improved | 408
granulation tissues | 408
transferred to a general ward | 408