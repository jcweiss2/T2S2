45 years old | 0
male | 0
admitted to hospital | 0
lizard bite | -48
severe pain | 0
marked swelling of the right leg | 0
decreased urine output | 0
conscious | 0
Glasgow coma scale E4V5M6 | 0
stable vitals | 0
respiratory distress | 24
respiratory rate 34-36/min | 24
oxygen saturation 85%-90% | 24
PaO2 64.1 mmHg | 24
FiO2 0.4 | 24
PCO2 22.7 mm Hg | 24
pH 7.29 | 24
bicarbonate 17.2 mmol/L | 24
BE -15.4 | 24
invasive mechanical ventilation | 24
total urine output 350 ml | 24
tea coloured urine | 24
extensive cellulitis | 24
marked oedema | 24
haemorrhagic bullae | 24
neutrophil leucocytosis | 48
intravascular haemolysis | 48
acute kidney injury | 48
injection tigecycline | 48
injection metronidazole | 48
normal saline infusion | 48
injection frusemide | 48
oliguric | 48
urinalysis | 48
reddish brown urine | 48
3+ protein | 48
pH 6 | 48
positive for blood | 48
20-25 red blood cells | 48
2-5 white blood cells | 48
rhabdomyolysis | 48
raised serum creatinine kinase | 48
raised serum myoglobin | 48
haemodialysis | 96
improved general condition | 192
weaned off ventilator | 144
decreasing trend of CK and myoglobin | 144
returned to normal on 13th day | 312
improved urine output | 360
nutrition with enteral renal formula | 360
oral renal diet | 360
shifted to ward | 432
discharged from hospital | 504