5 years old| 0
    male | 0
    emergency craniotomy | 0
    decompression of right parieto0occipital glioma | 0
    operated 3 months earlier | -4320
    worsening sensorium | -4320
    weakness of the left side | -4320
    Glasgow coma scale E2 V2 M3 | 0
    bilateral crackles | 0
    surgical emergency | 0
    ICU care | 0
    postoperative ventilator support | 0
    fasting state | 0
    blood grouping | 0
    cross matching | 0
    blood products arranged | 0
    sensorium deteriorating | 0
    no sedative premedication | 0
    ECG attached | 0
    SpO2 monitoring | 0
    noninvasive blood pressure monitoring | 0
    premedicated with fentanyl 40 mcg | 0
    induced with thiopental 100 mg | 0
    loss of eye lash reflex | 0
    bag0mask ventilation | 0
    vecuronium 2 mg | 0
    ventilated for 3 min | 0
    trachea intubated | 0
    endotracheal tube 5.5 mm ID | 0
    tube placement confirmed with capnography | 0
    tube secured at 15 cm | 0
    arterial line placed | 0
    left radial artery cannula 22-gauge | 0
    central line deferred | 0
    peripheral venous access | 0
    medial malleolar veins cannulas 18-gauge | 0
    Foley's catheter inserted | 0
    anesthesia maintained | 0
    oxygen and air mixture | 0
    isoflurane | 0
    vecuronium | 0
    propofol infusion | 0
    noncontrast computed tomography | 0
    midline shift | 0
    edema | 0
    arterial blood gas | 0
    mild hypocapnia 30–35 mm Hg | 0
    electrolyte correction | 0
    Mannitol 100 ml over 45 min | 0
    furosemide 10 mg | 0
    phenytoin | 0
    dexamethasone | 0
    antibiotics | 0
    surgery lasted 3 h | 0
    blood loss 400 ml | 0
    crystalloids replaced | 0
    packed red blood cells 200 ml transfused | 0
    preoperative GCS poor | 0
    ventilate patient | 0
    cerebral edema reduction | 0
    central venous access attempted | 0
    right subclavian approach | 0
    7 French Triple lumen B Braun central line | 0
    pilot puncture successful | 0
    guidewire insertion failed | 0
    ipsilateral internal jugular vein approach | 0
    guidewire advanced | 0
    no ECG rhythm changes | 0
    free blood flow from two ports | 0
    line secured with sutures | 0
    shifted to ICU | 0
    chest X-ray | 0
    central line malpositioned | 0
    no pneumothorax | 0
    line removed | 0
    peripheral venous access | 24
    Triple lumen B Braun Central Line inserted | 24
    left IJV approach | 24
    postoperative cardiovascular instability | 24
    sepsis | 24
    ventilatory support removed | 240
    shifted to surgical ward | 336
    