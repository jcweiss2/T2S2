26 years old | 0
female | 0
familial adenomatous polyposis | -672
prior proctocolectomy with J-pouch | -672
elective laparotomy with ileostomy reversal | 0
post-operative volvulus | 0
ischemic bowel with perforation | 0
emergent abdominal exploration | 0
small bowel resection | 0
drainage of abdominal and pelvic abscesses | 0
admitted to the intensive care unit | 0
hemodynamically unstable | 0
tachycardia to 190 beats per minute | 0
mean arterial pressure of 65 mm Hg | 0
central venous oxygen (SCVO2) value of 51% | 0
central venous pressure of 16 cmH2O | 0
positive fluid balance of 10 L | 0
vasopressin infusion | 0
epinephrine infusion | 0
norepinephrine infusion | 0
arterial blood gas analysis | 0
profound hypoxemia | 0
acidemia | 0
rising serum lactate level | 0
bilateral alveolar infiltrates | 0
atrial flutter with variable conduction | 0
Troponin I values mildly elevated | 0
transthoracic echocardiography | 0
TTS with regional wall motion abnormalities (RWMAs) | 0
akinet left ventricular apex | 0
compensatory hyperkinesis of the ventricle base | 0
moderate tricuspid valve regurgitation | 0
right ventricular systolic pressure of 60 mm Hg | 0
left ventricular ejection fraction (LVEF) approximately 15%–20% | 0
insertion of a left ventricular assist device | 0
left and right heart catheterization | 0
coronary angiogram | 0
insertion of a Swan-Ganz pulmonary arterial catheter | 0
Impella CP left ventricular assist device | 0
initial output set at 2.8 L/min | 0
no significant coronary obstructing lesions | 0
pulmonary arterial pressure | 0
mean pressure of 27 mm Hg | 0
wedge pressure of 25 mm Hg | 0
inhaled prostaglandins | 24
milrinone infusion | 24
improved oxygenation | 24
auto-anticoagulation | 24
thrombocytopenia | 24
systemic heparinization | 24
mild hematuria | 24
acute kidney injury | 48
device remained in situ without complications | 108
device removed | 108
hemodynamic improvement | 108
recovery of the ejection fraction to 40% | 108
discharged from the intensive care unit | 672
returned to almost full health | 1008