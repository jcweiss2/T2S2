70 years old | 0
male | 0
emergency esophageal diversion | -156
injury to the cervical esophagus | -156
spinal surgery | -156
gastric pull-up procedure | -132
postoperative anastomotic leakage | -132
endoscopy | -132
esophageal stent | -132
discharged | -114
local cervical infection | -102
sepsis | -102
admitted to hospital | 0
malnutrition | 0
systemic inflammation | 0
jugular and cervical phlegmon | 0
hemoglobin level of 6.7 g/dL | 0
white blood cell count of 6400 cells/μL | 0
platelet count of 210 × 103/μL | 0
creatinine level of 0.76 mg/dL | 0
albumin level of 2.8 g/dL | 0
chest computed tomography scan | 0
endoscopy | 0
dislodged esophageal stent | 0
esophageal perforation | 0
infected cavity | 0
esophageal stenosis | 0
stent removal | 0
endoscopic vacuum therapy | 12
EsoSponge system | 12
jugular and cervical phlegmon resolved | 168
repeated endoscopic balloon dilatation | 168
subtotal esophageal resection | 336
reconstruction using a free-jejunal graft interposition | 336
CT angiography | 336
partial sternotomy | 336
laparotomy | 336
jejunal segment harvested | 336
left carotid artery and left jugular vein used as recipient vessels | 336
graft implanted in an isoperistaltic position | 336
cervical anastomosis performed in an end-to-end fashion | 336
upper mediastinal gastro-jejunostomy performed in a side-to-side fashion | 336
upper sternum resected | 336
soft tissue defect covered with a sternocleidomastoid muscle flap | 336
abdominal reconstruction achieved by an end-to-end jejunojejunostomy | 336
postoperative course uneventful | 360
oral alimentation reestablished | 360
speech therapy | 360
anastomotic healing confirmed radiologically and endoscopically | 360
transferred to a rehabilitation clinic | 360
arterial hypertonus | -156
non-active smoking status | -156
ischemic stroke with incomplete senso-motoric hemiparesis | -156
thyroidectomy | -156
open prostatectomy due to prostate cancer | -156
family history not related to present illness | 0
personal history | 0