56 years old | 0
male | 0
intermittent headache | -72
fever | -72
transsphenoidal surgery | -2628
subtotal tumor resection for pituitary adenoma | -2628
gamma knife stereo-radiosurgery | -2628
gamma knife stereo-radiosurgery | -700
body temperature 38.2°C | 0
heart rate 85 bpm | 0
blood pressure 125/78 mm Hg | 0
respiratory rate 18 breaths/min | 0
doubtful neck resistance | 0
right pupil slightly larger | 0
asthenocoria | 0
oculomotor nerve injury | -2628
WBC count 10.12 × 10^9/L | 0
neutrophil ratio 59.9% | 0
CRP 12.9 mg/L | 0
blood glucose 6.63 mmol/L | 0
D-dimer 860 μg/L | 0
coagulation test | 0
serum pituitary hormone test | 0
ECG studies | 0
chest CT scan | 0
abdominal ultrasonography | 0
CT scan | 0
residual tumor in sellar region | 0
suspicious hemorrhage | 0
dehydration therapy | 0
hemostasis therapy | 0
progressive headache | 3
loss of vision in left eye | 3
loss of consciousness | 3
arrest of spontaneous heartbeat and breath | 3
CPR | 3
head CT scan | 3
MR and MRV | 3
inhomogeneous CSF signal | 3
mechanical ventilation | 3
intensive care | 3
endotracheal intubation | 3
lumbar puncture | 48
intracranial pressure 400 mm H2O | 48
yellow and thick CSF | 48
CSF cytology | 48
purulent meningitis | 48
septic shock | 48
daptomycin and linezolid and voriconazole | 48
aerobic and anaerobic cultures | 48
CSF culture | 48
antibiotic sensitivity test | 48
K pneumoniae | 48
meropenem and vancomycin | 72
lateral ventricular drainage | 72
bilateral ventricular irrigation | 72
cardiac arrest | 96
death | 96