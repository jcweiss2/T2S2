35 years old | 0  
    female | 0  
    acute lymphocytic leukemia (in remission since 1997) | 0  
    diabetes mellitus | 0  
    bipolar disorder | 0  
    recurrent urinary tract infections | 0  
    obesity | 0  
    gastric bypass surgery | 0  
    presented with altered mental status | 0  
    bedbound for 3 months | -2160  
    withdrawn | -2160  
    decreased appetite | -2160  
    poor nutrition | -2160  
    tachycardic (150 bpm) | 0  
    tachypneic (30-40 bpm) | 0  
    hypotensive (72/52 mm Hg) | 0  
    severe cachexia | 0  
    mottled bilateral upper extremities | 0  
    necrotic sacral decubitus ulcer | 0  
    sluggish bilateral pupils | 0  
    right-sided downward gaze preference | 0  
    roving eye movements | 0  
    pH 7.564 | 0  
    PCO2 23 mm Hg | 0  
    PO2 67 mm Hg | 0  
    lactic acid 5.3 mmol/L | 0  
    leukocytosis (19.2 K/UL) | 0  
    neutrophilic predominance | 0  
    sodium 137 mmol/L |$