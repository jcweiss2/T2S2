67 years old|0  
    female|0  
    admitted to the emergency department|0  
    abdominal pain|-72  
    bleeding diarrhoea|-72  
    nausea|-72  
    hypertension|0  
    type 2 diabetes mellitus|0  
    dyslipidemia|0  
    blood pressure 95/71 mmHg|0  
    temperature 36.3 °C|0  
    oxygen saturation 92%|0  
    diffuse abdominal pain without peritonitis|0  
    leukocytes 7.3 × 10³ μL|0  
    hemoglobin 12.6 g/dL|0  
    platelet count 96 × 10³ μL|0  
    serum creatinine 1.45 mg/dL|0  
    serum sodium 132 mmol/L|0  
    serum potassium 4.5 mmol/L|0  
    acute gastroenteritis|0  
    acute prerenal failure|0  
    treated with fluids|0  
    proton pump inhibitor|0  
    antiemetics|0  
    intravenous antibiotic therapy with ciprofloxacin|0  
    intravenous antibiotic therapy with metronidazole|0  
    stool culture sent|0  
    continued anuria|-24  
    unfavourable evolution on blood test|0  
    non-significant schistocytes count (< 1%)|0  
    abdominal CT scan|-48  
    proctitis (inflammatory/infectious)|0  
    cortical hypoperfusion of both kidneys|0  
    admitted to intensive care unit (ICU)|72  
    neurological failure with bradipsiquia|72  
    anuria|72  
    worsen blood test analysis|72  
    no hemodynamic instability|72  
    no respiratory failure|72  
    hemoglobin 11.2 g/dL|72  
    haptoglobin < 6.63 mg/dL|72  
    lactate dehydrogenase 1125 U/L|72  
    elevated schistocytes count on blood smear|72  
    negative direct antiglobulin test|72  
    microangiopathic haemolytic anemia|72  
    thrombocytopenia (post transfusion platelet count 59 × 10³ μL)|72  
    diagnosed with TMA|72  
    treated with urgent plasma exchange|72  
    methylprednisolone 1 mg/kg per day|72  
    uremia requiring haemodialysis|72  
    ADAMTS13 test result (55.9%)|96  
    daily plasma exchange sessions|72  
    possible severe atypical HUS|72  
    deterioration of neurological situation|72  
    persistence of anuric renal failure|72  
    low C3 complement levels|72  
    plasma exchange discontinued|96  
    verotoxin 2-secreting Escherichia Coli isolated|96  
    favourable clinical evolution|96  
    improvement of neurological symptoms after third day|144  
    transferred to ward|120  
    slower renal failure improvement|168  
    recovery of diuresis at second week|336  
    haemodialysis until 23rd day|552  
    renal biopsy confirming thrombotic microangiopathic involvement|552  
    anemia increasing slowly|168  
    no red-cell transfusion until sixth day|144  
    marked platelet decrease requiring transfusion|72  
    invasive techniques requiring platelet transfusion|72  
    endothelial congestion in renal biopsy|552  
    mesangial cellularity causing vascular occlusion|552  
    aneurysmal dilation of glomerular capillaries|552  
    polymorphonuclear and fragmented erythrocytes|552  
    thrombotic microangiopathic involvement in initial acute phase|552  
    treatment with plasma exchange started at 4 hours|72  
    ADAMTS13 levels received in 24 hours|96  
    TTP ruled out|96  
    atypical HUS considered|72  
    eculizumab evaluated|96  
    verotoxin 2-secreting Escherichia Coli confirmed|96  
    typical HUS diagnosed|96  
    plasma exchange stopped|96  
    eculizumab not used|96  
    Shiga-toxin-induced endothelial damage|0  
    bloody diarrhoea from verotoxin|0  
    supportive treatment|72  
    antibiotics controversial|72  
    plasma exchange no benefit|96  
    eculizumab uncertain role|96  
    neurological involvement|72  
    haemodialysis needed|72  
    complete renal recovery in four weeks|672  
    no financial support received|0  
    Institutional Ethics Committee approval|0  
    patient consent obtained|0  
    conflict of interest none|0  
    manuscript invited|0  
    critical care specialty|0  
    Spain origin|0  
    peer-review reports obtained|0  
    article in press|0  
    </s>

67 years old|0  
female|0  
admitted to the emergency department|0  
abdominal pain|-72  
bleeding diarrhoea|-72  
nausea|-72  
hypertension|0  
type 2 diabetes mellitus|0  
dyslipidemia|0  
blood pressure 95/71 mmHg|0  
temperature 36.3 °C|0  
oxygen saturation 92%|0  
diffuse abdominal pain without peritonitis|0  
leukocytes 7.3 × 10³ μL|0  
hemoglobin 12.6 g/dL|0  
platelet count 96 × 10³ μL|0  
serum creatinine 1.45 mg/dL|0  
serum sodium 132 mmol/L|0  
serum potassium 4.5 mmol/L|0  
acute gastroenteritis|0  
acute prerenal failure|0  
treated with fluids|0  
proton pump inhibitor|0  
antiemetics|0  
intravenous antibiotic therapy with ciprofloxacin|0  
intravenous antibiotic therapy with metronidazole|0  
stool culture sent|0  
continued anuria|-24  
unfavourable evolution on blood test|0  
non-significant schistocytes count (< 1%)|0  
abdominal CT scan|-48  
proctitis (inflammatory/infectious)|0  
cortical hypoperfusion of both kidneys|0  
admitted to intensive care unit (ICU)|72  
neurological failure with bradipsiquia|72  
anuria|72  
worsen blood test analysis|72  
no hemodynamic instability|72  
no respiratory failure|72  
hemoglobin 11.2 g/dL|72  
haptoglobin < 6.63 mg/dL|72  
lactate dehydrogenase 1125 U/L|72  
elevated schistocytes count on blood smear|72  
negative direct antiglobulin test|72  
microangiopathic haemolytic anemia|72  
thrombocytopenia (post transfusion platelet count 59 × 10³ μL)|72  
diagnosed with TMA|72  
treated with urgent plasma exchange|72  
methylprednisolone 1 mg/kg per day|72  
uremia requiring haemodialysis|72  
ADAMTS13 test result (55.9%)|96  
daily plasma exchange sessions|72  
possible severe atypical HUS|72  
deterioration of neurological situation|72  
persistence of anuric renal failure|72  
low C3 complement levels|72  
plasma exchange discontinued|96  
verotoxin 2-secreting Escherichia Coli isolated|96  
favourable clinical evolution|96  
improvement of neurological symptoms after third day|144  
transferred to ward|120  
slower renal failure improvement|168  
recovery of diuresis at second week|336  
haemodialysis until 23rd day|552  
renal biopsy confirming thrombotic microangiopathic involvement|552  
anemia increasing slowly|168  
no red-cell transfusion until sixth day|144  
marked platelet decrease requiring transfusion|72  
invasive techniques requiring platelet transfusion|72  
endothelial congestion in renal biopsy|552  
mesangial cellularity causing vascular occlusion|552  
aneurysmal dilation of glomerular capillaries|552  
polymorphonuclear and fragmented erythrocytes|552  
thrombotic microangiopathic involvement in initial acute phase|552  
treatment with plasma exchange started at 4 hours|72  
ADAMTS13 levels received in 24 hours|96  
TTP ruled out|96  
atypical HUS considered|72  
eculizumab evaluated|96  
verotoxin 2-secreting Escherichia Coli confirmed|96  
typical HUS diagnosed|96  
plasma exchange stopped|96  
eculizumab not used|96  
Shiga-toxin-induced endothelial damage|0  
bloody diarrhoea from verotoxin|0  
supportive treatment|72  
antibiotics controversial|72  
plasma exchange no benefit|96  
eculizumab uncertain role|96  
neurological involvement|72  
haemodialysis needed|72  
complete renal recovery in four weeks|672  
no financial support received|0  
Institutional Ethics Committee approval|0  
patient consent obtained|0  
conflict of interest none|0  
manuscript invited|0  
critical care specialty|0  
Spain origin|0  
peer-review reports obtained|0  
article in press|0  
