51 years old | 0
    male | 0
    asthma | -672
    unconscious | -16
    taken to local clinic | -16
    taken to regional hospital | -16
    swallowed agricultural pesticide (organophosphate) | -16
    Atropine Challenge test (negative) | -16
    intubated due to loss of consciousness (GCS 8) | -16
    sent to poison centers | -16
    blood pressure 65/40 mmHg | -16
    metabolic acidosis | -16
    consultation with subspecialized center (clinical toxicology) | -16
    possibility of aluminum phosphide poisoning | -16
    treated with normal saline | -16
    norepinephrine infusion | -16
    bicarbonate | -16
    hydrocortisone | -16
    loading dose of NAC | -16
    clarified ingestion of 1 liter hexaflumuron 10% | -16
    no evidence of pills or other poisons | -16
    transferred to Imam Reza Toxicology Center | 0
    GCS 5 on admission | 0
    BP 78/36 mmHg | 0
    pulse rate 80 beats/min | 0
    axillary temperature 37.2°C | 0
    respiratory rate 22 cycles/min | 0
    intubated | 0
    mechanically ventilated (SIMV) | 0
    pupils normal | 0
    cherry-colored skin on lower limbs and abdomen | 0
    blood glucose 204 mg/dL | 0
    fluid therapy | 0
    cardiac monitoring | 0
    ventilated | 0
    reduced blood pressure | 0
    no manifestations of organophosphate poisoning | 0
    aluminum phosphide poisoning treatment | 0
    administered norepinephrine | 0
    hydrocortisone 200 mg IV | 0
    NAC 140 mg/kg IV | 0
    carboxyhemoglobin level tested | 0
    urine paraquat test | 0
    serum cholinesterase levels | 0
    red blood cell cholinesterase levels | 0
    urine immunoassay positive for tricyclic antidepressant | 0
    no blocking cardiac sodium channel on ECG | 0
    QTc 0.56 | 0
    magnesium sulfate 2 g | 0
    magnesium sulfate repeated every 8 hours | 0
    echocardiogram normal wall motion (EF 55%) | 0
    transferred to ICU 3 hours after admission | 3
    blood pressure 80/50 at 4:15 PM | 3
    re-administered 1 liter normal saline | 3
    VBG values analyzed | 3
    suspicion of aluminum phosphide poisoning | 3
    100 mEq bicarbonate administered | 3
    continued bicarbonate infusion | 3
    potassium supplementation | 3
    white blood cell count 21.81 *1000/µL | 0
    hemoglobin 15.1 g/dL | 0
    hematocrit 44.5% | 0
    platelet 434 *1000/µL | 0
    neutrophil 53% | 0
    lymphocyte 44% | 0
    PT 15.4 sec | 0
    INR 1.49 | 0
    PTT 30 sec | 0
    pH 7.039 | 0
    PCO2 43.8 mmHg | 0
    HCO3 11.8 mEq/L | 0
    base excess -19.0 mmol/L | 0
    PO2 115.5 mmHg | 0
    O2 saturation 95.5% | 0
    sodium 138 mg/dL | 0
    potassium 3.3 mg/dL | 0
    chloride 114 mg/dL | 0
    calcium 8.7 mg/dL | 0
    phosphorus 2.2 mg/dL | 0
    magnesium 2.7 mg/dL | 0
    urea 28 mg/dL | 0
    creatinine 2.1 mg/dL | 0
    blood sugar 247 mg/dL | 0
    lactate dehydrogenase 622 U/L | 0
    creatine phosphokinase 444 U/L | 0
    AST 40 U/L | 0
    ALT 23 U/L | 0
    alkaline phosphatase 181 U/L | 0
    total bilirubin 0.88 mg/dL | 0
    direct bilirubin 0.24 mg/dL | 0
    troponin I 8.5 | 0
    NT pro BNP 1142 Pg/ML | 0
    procalcitonin 0.92 ng/ml | 0
    norepinephrine infusion discontinued (30 hours after admission) | 30
    decreased QTc intervals | 30
    magnesium sulfate discontinued | 30
    serum creatinine 2.6 mg/dL | 30
    low urinary volume | 30
    furosemide administered | 30
    urine output appropriate | 30
    fluid therapy continued | 30
    bicarbonate continued | 30
    metabolic acidosis improvement | 54
    bicarbonate discontinued | 54
    not ready for ventilator withdrawal | 54
    pulmonary edema | 54
    morphine administered | 54
    furosemide administered | 54
    echocardiogram normal | 54
    pneumonia (pulmonary x-ray) | 54
    antibiotic treatment started | 54
    broncho-vascular markings increased | 54
    para-cardiac opacity | 54
    patchy opacity in both lungs | 54
    uniform opacity in right lung | 54
    blood culture performed | 54
    urine culture performed | 54
    urine culture positive for E. coli | 54
    blood culture negative | 54
    fever developed | 54
    fever treatment | 54
    bradycardia | 96
    hypotension | 96
    cardiac arrest | 96
    cardiopulmonary resuscitation | 96
    death | 96
    <|eot_id|>
    51 years old | 0
male | 0
asthma | -672
unconscious | -16
taken to local clinic | -16
taken to regional hospital | -16
swallowed agricultural pesticide (organophosphate) | -16
Atropine Challenge test (negative) | -16
intubated due to loss of consciousness (GCS 8) | -16
sent to poison centers | -16
blood pressure 65/40 mmHg | -16
metabolic acidosis | -16
consultation with subspecialized center (clinical toxicology) | -16
possibility of aluminum phosphide poisoning | -16
treated with normal saline | -16
norepinephrine infusion | -16
bicarbonate | -16
hydrocortisone | -16
loading dose of NAC | -16
clarified ingestion of 1 liter hexaflumuron 10% | -16
no evidence of pills or other poisons | -16
transferred to Imam Reza Toxicology Center | 0
GCS 5 on admission | 0
BP 78/36 mmHg | 0
pulse rate 80 beats/min |0
axillary temperature 37.2°C | 0
respiratory rate 22 cycles/min | 0
intubated | 0
mechanically ventilated (SIMV) | 0
pupils normal | 0
cherry-colored skin on lower limbs and abdomen | 0
blood glucose 204 mg/dL | 0
fluid therapy | 0
cardiac monitoring | 0
ventilated | 0
reduced blood pressure | 0
no manifestations of organophosphate poisoning | 0
aluminum phosphide poisoning treatment | 0
administered norepinephrine | 0
hydrocortisone 200 mg IV | 0
NAC 140 mg/kg IV | 0
carboxyhemoglobin level tested | 0
urine paraquat test | 0
serum cholinesterase levels | 0
red blood cell cholinesterase levels | 0
urine immunoassay positive for tricyclic antidepressant | 0
no blocking cardiac sodium channel on ECG | 0
QTc 0.56 | 0
magnesium sulfate 2 g | 0
magnesium sulfate repeated every 8 hours | 0
echocardiogram normal wall motion (EF 55%) | 0
transferred to ICU 3 hours after admission | 3
blood pressure 80/50 at 4:15 PM | 3
re-administered 1 liter normal saline | 3
VBG values analyzed | 3
suspicion of aluminum phosphide poisoning | 3
100 mEq bicarbonate administered | 3
continued bicarbonate infusion | 3
potassium supplementation | 3
white blood cell count 21.81 *1000/µL | 0
hemoglobin 15.1 g/dL | 0
hematocrit 44.5% | 0
platelet 434 *1000/µL | 0
neutrophil 53% | 0
lymphocyte 44% | 0
PT 15.4 sec | 0
INR 1.49 | 0
PTT 30 sec | 0
pH 7.039 | 0
PCO2 43.8 mmHg | 0
HCO3 11.8 mEq/L | 0
base excess -19.0 mmol/L | 0
PO2 115.5 mmHg | 0
O2 saturation 95.5% | 0
sodium 138 mg/dL | 0
potassium 3.3 mg/dL | 0
chloride 114 mg/dL | 0
calcium 8.7 mg/dL | 0
phosphorus 2.2 mg/dL | 0
magnesium 2.7 mg/dL | 0
urea 28 mg/dL | 0
creatinine 2.1 mg/dL | 0
blood sugar 247 mg/dL | 0
lactate dehydrogenase 622 U/L | 0
creatine phosphokinase 444 U/L | 0
AST 40 U/L | 0
ALT 23 U/L | 0
alkaline phosphatase 181 U/L | 0
total bilirubin 0.88 mg/dL | 0
direct bilirubin 0.24 mg/dL | 0
troponin I 8.5 | 0
NT pro BNP 1142 Pg/ML | 0
procalcitonin 0.92 ng/ml | 0
norepinephrine infusion discontinued (30 hours after admission) | 30
decreased QTc intervals | 30
magnesium sulfate discontinued | 30
serum creatinine 2.6 mg/dL | 30
low urinary volume | 30
furosemide administered | 30
urine output appropriate | 30
fluid therapy continued | 30
bicarbonate continued | 30
metabolic acidosis improvement | 54
bicarbonate discontinued | 54
not ready for ventilator withdrawal | 54
pulmonary edema | 54
morphine administered | 54
furosemide administered | 54
echocardiogram normal | 54
pneumonia (pulmonary x-ray) | 54
antibiotic treatment started | 54
broncho-vascular markings increased | 54
para-cardiac opacity | 54
patchy opacity in both lungs | 54
uniform opacity in right lung | 54
blood culture performed | 54
urine culture performed | 54
urine culture positive for E. coli | 54
blood culture negative | 54
fever developed | 54
fever treatment | 54
bradycardia | 96
hypotension | 96
cardiac arrest | 96
cardiopulmonary resuscitation | 96
death | 96