55 years old | 0
male | 0
Caucasian | 0
admitted to hospital | 0
common cold | -168
myalgia | -168
fatigue | -168
headaches | -168
pleuritic chest pain | -168
breathlessness on exertion | -168
mild asthma | 0
Beclomethasone 100 µg, 2 puffs bd | 0
salbutamol 100 µg, 2 puffs prn | 0
ex-smoker | 0
25-pack years | 0
body mass index 24.6 kg/m2 | 0
blood pressure 130/80 mmHg | 0
pulse 110 bpm | 0
temperature 38.2°C | 0
decreased air entry on the right lung | 0
coarse crackles | 0
normal heart sounds | 0
no murmurs | 0
sinus tachycardia | 0
PR interval 124 ms | 0
QRS duration 99 ms | 0
corrected QT interval 382 ms | 0
no ST-T wave abnormalities | 0
serum creatinine 85 umol/L | 0
alanine aminotransferase 216 IU/L | 0
potassium level 5.4 mmoL/mL | 0
magnesium 1.2 | 0
corrected calcium 2.26 | 0
sodium 138 | 0
C-reactive protein 184 mg/L | 0
haemoglobin 86 g/L | 0
normocytic, normochromic | 0
platelets 670 × 109/L | 0
WBC 18 × 109/L | 0
neutrophilia | 0
international normalised ratio 1.4 | 0
activated partial thromboplastin time 27.2 s | 0
right sided consolidation | 0
Pseudomonas aeruginosa | 0
oxygen | 0
intravenous fluids | 0
antibiotics | 0
meropenem | 0
clarithromycin | 0
central chest pain | -96
inferior ST elevation myocardial infarction | -96
drug eluting stent to left circumflex coronary artery | -96
atrial fibrillation | -96
ventricular bigeminy | -96
dual antiplatelet therapy | -96
aspirin | -96
ticagrelor | -96
respiratory deterioration | -72
intubation | -72
invasive ventilation | -72
veno-venous extracorporeal membrane oxygenation | -72
atrial fibrillation with ventricular rate 140–150 bpm | -60
ventricular ectopy | -60
run of ventricular tachycardia | -60
increasing noradrenaline requirement | -60
mean arterial pressure 59 mmHg | -60
amiodarone loading | -60
repeated angiogram | -48
patent LCx stent | -48
left anterior descending disease | -48
treated with 2 DES | -48
atrial fibrillation with fast ventricular rate | -36
esmolol | -36
bradycardia | -36
VF arrest | -36
Torsade de Pointes | -36
corrected QT interval 550 ms | -36
CPR | -36
direct current cardioversion | -36
return of spontaneous circulation | -36
post arrest ECG | -36
persistent VE | -24
AF | -24
bradycardic episodes | -24
increase in noradrenaline requirement | -24
atrial pacemaker | -12
AAI 90 bpm | -12
cessation of VE | 0
cessation of AF | 0
reduction in noradrenaline requirement | 0
decannulated from ECMO | 12
insertion of secondary-prevention implantable cardioverter defibrillator | 24
repatriated to local ICU | 48
died of sepsis | 72