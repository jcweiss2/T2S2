46 years old | 0
male | 0
admitted to ICU | 0
severe chronic obstructive pulmonary disease (COPD) | 0
bronchial asthma | 0
acute proptosis of both eyes | 0
globe luxation | 0
retracted lids | 0
history of similar episode in the past | -8760
previous episodes over past 4–5 years | -8760
wheezing episodes | -8760
exacerbations of COPD | -8760
bilateral pseudophakia | 0
normal pupil | 0
normal fundus | 0
axial length in both eyes was 23.8 mm | 0
computed tomography (CT) scan of orbit | 0
no orbital mass | 0
proptosed eye with a stretched optic nerve | 0
orbit volume and globe volume appeared normal | 0
repeated episodes of globe luxation | 2
repeated episodes of globe luxation | 4
repeated episodes of globe luxation | 6
bilateral temporary tarsorrhaphy | 12
respiratory paralysis | 48
septicemia | 48
expired | 72
globe luxation reduced | 0
globe luxation reduced | 2
globe luxation reduced | 4
globe luxation reduced | 6
Valsalva maneuver | -8760
lid manipulation | -8760
trauma | -8760
general anesthesia | -8760
contact lens insertion | -8760
histiocytosis X | -8760
Engelmann's disease | -8760
thyroid eye disease | -8760
floppy eyelid syndrome | -8760
shallow orbit | -8760
lateral tarsorrhaphy | 12
pentagonal wedge eyelid resection | -8760
advancement of orbital wall | -8760