24 years old | 0
    female | 0
    presented to the emergency department | 0
    severe headache | -72
    projectile vomiting | -72
    no history of fever | 0
    no history of convulsions | 0
    no history of focal neurological deficit | 0
    treated outside symptomatically | -72
    no relief | -72
    provisionally diagnosed with metabolic encephalopathy | 0
    symptomatic treatment | 0
    transferred to intensive care unit | 24
    deteriorated further | 24
    altered sensorium (GCS-9) | 24
    high-grade fever | 24
    chills | 24
    dyselectrolytemia (serum potassium – 3.7 mEq/L) | 24
    low serum phosphate (1.57 mg/dL) | 24
    neutrophilic leukocytosis (TLC – 24,170/μl, neutrophils – 91%) | 24
    cerebrospinal fluid sent for evaluation | 24
    empirically treated with ceftriaxone | 24
    Gram stain of CSF deposit revealed polymorphs and lymphocytes | 24
    Gram-positive bacilli in CSF | 24
    culture of CSF grew Listeria monocytogenes | 24
    conventional identification methods | 24
    automated methods (VITEK-2) | 24
    blood culture taken at admission grew Gram-positive bacilli | 0
    ignored as diphtheroids | 0
    reevaluation recognized as L. monocytogenes | 24
    similar sensitivity pattern | 24
    switched to meropenem | 48
    other corrective measures | 48
    clinical improvement | 48
    microbiological improvement | 48
    CSF biochemistry: raised protein (91 mg/dL) | 24
    CSF biochemistry: decreased glucose (6 mg/dL) | 24
    CSF biochemistry: normal ADA | 24
    CSF cytology: high cell count (1080/cm) | 24
    CSF cytology: 60% neutrophils | 24
    CSF cytology: 40% lymphocytes | 24
    Gram-positive bacilli in blood culture | 0
    meningitis due to L. monocytogenes | 24
    no preexisting illness | 0
    no prolonged medication | 0
    lower incidence of meningeal signs | 24
    dyselectrolytemia | 24
    inherent resistance to cephalosporin | 24
    inherent resistance to vancomycin | 24
    microbiological diagnosis | 24
    identification challenging due to diphtheroids appearance | 24
    identification challenging due to diplococci appearance | 24
    contamination risk | 24
    listerial infection in young healthy adults | 24
    careful microbiological identification | 24
    proper diagnosis | 24
    treatment | 24
    declaration of patient consent | 0
    no financial support | 0
    no conflicts of interest | 0