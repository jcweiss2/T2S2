10-year-old | 0
    boy | 0
    born pre-term | 0
    gestational age of 33 weeks and 2 days | 0
    developmental delays in growth | 0
    developmental delays in motor function | 0
    first visited our center for evaluation of short stature | -35040
    clinical diagnosis with Russell–Silver syndrome | -35040
    proteinuria | -35040
    hypoalbuminemia | -35040
    high-dose steroid | -35040
    calcineurin inhibitor | -35040
    deteriorated renal function | -35040
    right renal vein thrombosis | -17544
    pulmonary embolism | -17544
    treated with anticoagulants | -17544
    persistent pulmonary hypertension | -17544
    managed with sildenafil | -17544
    underwent living donor kidney transplantation | -8760
    immunosuppression using prednisolone | -8760
    mycophenolate mofetil (MMF) | -8760
    tacrolimus | -8760
    discontinued MMF | -8760 + 70 days (70 days after transplantation)
    steroid was tapered | -8760 + 70 days
    tacrolimus continued with blood levels maintained at approximately 10 ng/mL | -8760 + 70 days
    developed pneumocystis pneumonia | -8760 + 70 days + 3 months (approx 3 months after transplantation)
    necessitated mechanical ventilation | -8760 + 70 days + 3 months
    treated with intravenous sulfamethoxazole/trimethoprim for 14 days | -8760 + 70 days + 3 months
    steroid increased from 2.5 mg to 20 mg prednisolone | -8760 + 70 days + 3 months
    continued at same dose after discharge | -8760 + 70 days + 3 months + 14 days (approx)
    presented with dysuria | 135 days post-transplantation (0 at admission)
    presented with gross hematuria | 135 days post-transplantation (0 at admission)
    BUN 24 mg/dL | 0
    Cr 0.56 mg/dL | 0
    CRP 0.42 mg/dL | 0
    RBC count > 100/HPF | 0
    WBC count > 100/HPF | 0
    urine culture for bacteria negative | 0
    BK virus negative | 0
    urine JC virus PCR positive | 0
    urine adenovirus culture positive (1–9 cells/HPF) | 0
    diagnosed with hemorrhagic cystitis | 0
    managed with hydration | 0
    managed with pain control | 0
    dysuria persisted | +168 (1 week after admission)
    hematuria persisted | +168
    RBC count > 100/HPF | +168
    WBC count 1 to 4/HPF | +168
    immunosuppression maintained | +168
    visited emergency room with fever | +504 (3 weeks after admission)
    general weakness | +504
    chest tightness | +504
    mild cough | +504
    persistent dysuria | +504
    persistent hematuria | +504
    BUN 175 mg/dL | +504
    Cr 8.29 mg/dL | +504
    CRP 30.23 mg/dL | +504
    emergent hemodialysis | +504
    empirically treated with piperacillin/tazobactam | +504
    sputum culture negative | +504
    blood culture negative | +504
    urine culture negative | +504
    adenovirus real-time PCR of sputum positive | +504
    blood CMV antigen positive | +504
    presumed disseminated adenovirus infection | +504
    treated with immunosuppression reduction | +504
    treated with ganciclovir | +504
    renal allograft biopsy showing diffuse necrotizing granulomatous tubulointerstitial nephritis | +504
    CD3 staining negative | +504
    C4d staining negative | +504
    positive JC virus PCR | +504
    serum CMV PCR positive | +504
    treated with ganciclovir targeting CMV | +504
    antibiotic therapy with renal impairment dose for CMV infection | +504
    granulocyte colony-stimulating factor | +504
    immunoglobulin | +504
    transfusion | +504
    hemodialysis | +504
    high inflammatory marker | +504
    persistent fever | +504
    initiated cidofovir treatment | +792 (167th day post-transplantation)
    given cidofovir 1 mg/kg/day 3 times/week without probenecid | +792
    changed regimen to 2 mg/kg every 2 weeks | +792 + ... (after 4 doses)
    serum adenovirus PCR positive | +792 + ...
    cerebrospinal fluid adenovirus PCR positive | +792 + ...
    renal function not recovered | +792 + ...
    generalized tonic-clonic seizure | +792 + ...
    treated with vancomycin | +792 + ...
    treated with meropenem | +792 + ...
    treated with acyclovir | +792 + ...
    anemia | +792 + ...
    leukopenia | +792 + ...
    thrombocytopenia | +792 + ...
    mechanical ventilation | +792 + ...
    continuous renal replacement therapy | +792 + ...
    died | +5160 (215th day post-transplantation)