88 years old | 0
female | 0
transferred to hospital with right hip pain | -432
fall while walking using a walker | -432
history of hypertension | 0
history of dementia | 0
conservative observation at home | -432
no improvement in hip pain | -432
visited another hospital | -432
diagnosed with intertrochanteric fracture | -432
planned surgical treatment | -432
preoperative evaluation diagnosed with COVID-19 | -432
transferred to isolation ward | -432
blood pressure drop to 94/39 mmHg | -432
urinary tract infection | -432
sepsis | -432
ischemic colitis | -432
transferred to ICU | -432
delayed planned surgery | -432
treatment for ischemic colitis | -432
treatment for septic shock | -432
transferred to current hospital | 0
surgical treatment 18 days after injury | 0
preoperative laboratory findings | 0
hemoglobin 9.0 g/dl | 0
platelet 169,000 µl | 0
serum albumin 3.28 g/dl | 0
C-reactive protein 2.7 mg/dl | 0
sodium 139 mEq/L | 0
arterial blood gas analysis | 0
pH 7.55 | 0
pCO2 37 mmHg | 0
PO2 63 mmHg | 0
HCO3- 32.1 mmol/L | 0
SaO2 94.1% | 0
prothrombin time 14.8 s | 0
international normalized ratio 1.21 | 0
activated partial thromboplastin time 35.3 s | 0
D-dimer 18.94 µg/ml | 0
chest CT showing diffuse PTE | 0
consolidation in right lower lobe | 0
ground glass opacity in both lower lobes | 0
small amount of right pleural effusion | 0
left rib fractures | 0
abdominopelvic CT showing DVT | 0
transthoracic echocardiography findings | 0
65% ejection fraction | 0
mild aortic stenosis | 0
thickened and calcified mitral valve | 0
trivial mitral regurgitation | 0
visible echogenic material in left atrium | 0
electrocardiography showed no atrial fibrillation | 0
cardiology consultation recommended delayed surgery 2-3 days after heparinization | 0
insertion of IVC filter | 0
admitted to operating room for right hip hemiarthroplasty | 0
preoperative vital signs | 0
BP 165/78 mmHg | 0
heart rate 72 beats/min | 0
body temperature 36.5℃ | 0
respiratory rate 20/min | 0
oxygen saturation 91% | 0
continuous radial arterial pressure monitoring | 0
TOF monitoring | 0
BIS monitoring | 0
anesthesia induced | 0
remimazolam administration | 0
rocuronium administration | 0
tracheal intubation performed | 0
anesthesia maintained | 0
remifentanil administration | 0
ECMO preparation | 0
introducer sheath inserted | 0
TEE probe inserted | 0
no thrombus observed in left atrium | 0
mean arterial pressure maintained over 70 mmHg | 0
ephedrine bolus administered | 0
fluid administered 1,400 ml plasmalyte | 0
bleeding 300 ml | 0
urine output 90 ml | 0
total anesthetic time 190 min | 0
total operating time 170 min | 0
flumazenil administration | 0
pyridostigmine administration | 0
glycopyrrolate administration | 0
tracheal extubation | 0
transferred to ICU | 0
ECMO sheaths removed | 48
transferred to general ward | 48
IVC filter removed | 192
discharged | 192
