27 years old | 0
female | 0
bilateral liposuction of the thighs | -240
liposuction of the abdomen | -240
bilateral fat grafting to the breasts | -240
fever | -168
bilateral breast pain | -168
paracetamol | -168
no antibiotic therapy | -168
symptoms progressed | -144
erythema | -144
swelling | -144
pain | -144
septic shock | 0
hypotension | 0
redness | 0
aggressive fluid resuscitation | 0
inotropes | 0
empirical intravenous penicillin G | 0
clindamycin | 0
ceftazidime | 0
computed tomography scans | 0
ill-defined masses | 0
sub-glandular planes | 0
air-fluid level | 0
surgery | 0
debridement | 0
foul-smelling fluid | 0
necrotic fat | 0
evacuation | 0
repeat debridement | 24
unhealthy tissue removed | 24
third debridement | 48
involvement of the left sternocleidomastoid muscle | 48
sepsis improved | 48
adequate debridement | 48
washout | 48
antibiotics | 48
supportive therapy | 48
bacterial cultures | 48
Proteus mirabilis | 48
Enterobacter aerogenes | 48
Enterococcus faecalis | 48
Bacteroides fragilis | 48
antibiotic therapy adjusted | 48
piperacillin-tazobactam | 48
further debridement operations | 72
wounds closed | 120
skin graft | 120
hypertrophic scars | 4320
follow-up | 4320