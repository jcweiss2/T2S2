51 years old | 0
male | 0
Caucasian | 0
admitted to the hospital | 0
dyspnoea | 0
peripheral pitting oedema | 0
orthopnoea | 0
paroxysmal nocturnal dyspnoea | 0
exercise tolerance limited to 40-50 m | 0
no chest pain | 0
no abdominal pain | 0
no palpitations | 0
no syncope | 0
no history of smoking | 0
no excessive alcohol consumption | 0
no drug use | 0
urosepsis | -7872
pyelonephritis | -7872
haemofiltration | -7872
CT scan | -7872
no cardiac changes | -7872
cardiomegaly | -768
moderate pericardial effusion | -768
diffuse mid-wall myocardial calcification | -768
transthoracic echocardiogram | -736
mildly dilated left ventricular | -736
moderate systolic dysfunction | -736
cerebrovascular event | -168
large LV apical thrombus | -168
anticoagulation | -168
bilateral below-knee pitting oedema | 0
respiratory distress | 0
heart rate 80 beats/min | 0
blood pressure 140/90 mmHg | 0
respiratory rate 18 breaths/minute | 0
SpO2 98% on room air | 0
temperature 37.0°C | 0
non-displaced apex beat | 0
no palpable thrills or right ventricular heave | 0
S1 and S2 heart sounds | 0
no added sounds, murmurs, or lung crepitations | 0
electrocardiogram | 0
left atrial enlargement | 0
pathological inferior Q waves | 0
no acute T wave or ST segment changes | 0
cardiac CT | 0
mild coronary artery disease | 0
no significant stenosis | 0
diffuse LV mid-wall myocardial calcification | 0
LVEF 20% | 0
valsartan/sacubitril | 0
spironolactone | 0
frusemide | 0
atorvastatin | 0
bisoprolol | 0
warfarin | 0
cardiac magnetic resonance imaging | 264
LVEF 34% | 264
diffuse LV mid-myocardial late gadolinium enhancement | 264
prophylactic implantable cardioverter-defibrillator | 552
New York Heart Association class II functional status | 552
non-ischaemic cardiomyopathy | 0
septic myocardial calcification | -7872
dystrophic calcification | -7872
metastatic calcification | -7872
catecholamine excess | -7872
nitric oxide | -7872
inducible nitric oxide synthase | -7872
microvascular ischaemia | -7872
scar-related arrhythmia | 0
ventricular systolic dysfunction | 0
ventricular arrhythmias | 0
atrioventricular conduction disorders | 0