77 years old | 0
male | 0
admitted to hospital | 0
anorexia | 0
deranged liver enzymes | 0
no significant past medical history | 0
no significant risk factors for liver disease | 0
does not take regular medications | 0
denied abdominal pain | 0
denied altered bowel habits | 0
afebrile | 0
hemodynamically stable | 0
unremarkable abdominal examination | 0
cholestatic liver enzymes | 0
elevated alkaline phosphatase | 0
elevated gamma-glutamyl transferase | 0
elevated total bilirubin | 0
raised white blood cell count | 0
raised neutrophil count | 0
abdominal ultrasound | 0
no visible gallstones | 0
became febrile | 336
worsening ALP and GGT | 336
Escherichia Coli bacteraemia | 336
Klebsiella pneumoniae bacteraemia | 336
diagnostic computed tomography scan | 336
hypodense focal liver lesions | 336
multiple thrombosed portal vein branches | 336
pneumobilia in the liver’s left lobe | 336
infra-renal abdominal aortic aneurysm | 336
commenced on Piperacillin–Tazobactam | 336
commenced on Rivaroxaban | 336
initially responded well to medical therapy | 336
large volume hematemesis | 504
clinically unstable | 504
repeat CT abdomen | 504
interval increase in the size of the infra-renal AAA | 504
Rivaroxaban ceased | 504
urgent gastroscopy | 504
large blood clots in the gastric fundus and body | 504
pulsatile lesion at the second part of the duodenum | 504
emergency endovascular aneurysm repair | 504
admitted to the intensive care unit | 504
complained of acute right lower limb pain and swelling | 624
Doppler ultrasound | 624
CT abdomen angiogram | 624
extensive deep vein thrombosis | 624
commenced an intravenous heparin infusion | 624
experienced a second episode of hematemesis | 720
third gastroscopy | 720
bleeding duodenal fistula at the D2/3 junction | 720
communicating with the gallbladder | 720
cholecystoduodenal fistula | 720
second laparotomy | 720
fistula between the gallbladder to the lateral wall of the duodenum | 720
several stones and sludge in a contracted gallbladder | 720
6 mm stone in the ampulla | 720
fistula and the adjacent duodenal wall were repaired | 720
cholecystectomy performed | 720
further hematemesis | 744
third laparotomy | 744
deep ulcer in D3 | 744
another aortoenteric fistula with D3 | 744
aneurysm sac bleeding into the duodenum | 744
iliolumbar arteries and inferior mesenteric artery closed | 744
survived the surgeries | 744
admitted into ICU | 744
later discharged from hospital | 744
re-admitted 3 weeks later | 1104
passed away from an unrelated event | 1104