66 years old | 0
male | 0
admitted to the hospital | 0
rash | -48
erythemato-violaceous macules | -48
papules | -48
purpuric elements | -48
itch | -48
postblister erosions on the oral and nasal mucosa | -48
genital erosions | -48
deep fissures | -48
haematic crusts on the lips | -48
painful burning sensations | -48
prodromal flu-like symptoms | -48
fever | -48
fatigue | -48
malaise | -48
diabetes mellitus type II | 0
insulin treatment | 0
chronic kidney disease stage 5 | 0
chronic hemodialysis | 0
obstructive nephropathy | 0
right nephrostomy | 0
secondary renal hypertension | 0
mixed decompensated toxic cirrhosis | 0
alcohol intake | 0
hepatic encephalopathy | 0
insulin 10 UI b.i.d. | 0
amlodipine 5 mg q.d. | 0
carbamazepine 100 mg q.d. | 0
hospitalized for hemodialysis | -48
slightly itchy erythemato-papulous rash on the face, hands, feet | -48
extension of the rash | -24
appearance of purpuric elements | -24
tendency to spread | -24
appearance of flaccid blisters | 0
eruption of blisters | 0
large areas of denudation | 0
preliminary diagnosis of drug-induced allergic vasculitis | 0
transfer to the Department of Dermatology | 0
malaise at admission | 0
itchy rash | 0
erythemato-violaceous macules | 0
purpuric macules | 0
papules | 0
patches | 0
dissemination on the trunk, upper and lower limbs, cephalic extremities | 0
flaccid blisters | 0
erosions | 0
denudation over 10% of the skin | 0
oral mucosal erosions | 0
nasal mucosal erosions | 0
deep fissures | 0
haematic crusts | 0
genital mucosal erosions | 0
yellow-white exudates | 0
balano-preputial folding | 0
high blood pressure (160/120 mmHg) | 0
increased abdominal volume due to ascites | 0
collateral venous circulation on the abdominal wall | 0
absence of neurological manifestations | 0
marked anemia | 0
leukocytosis | 0
neutrophilia | 0
thrombocytopenia | 0
inflammatory syndrome | 0
elevated ASLO titer | 0
elevated IgE | 0
nitrogen retention syndrome | 0
elevated blood sugar levels | 0
hydro-electrolyte imbalance | 0
hypokalemia | 0
low RA | 0
abnormal liver function | 0
reversing albumin/globulin rate | 0
normal serum total proteins | 0
normal INR | 0
bacterial supra-infection with Klebsiella pneumoniae | 0
multi-resistant to antibiotics | 0
sensitive to colistin | 0
sensitive to amikacin | 0
sensitive to ertapenem | 0
sensitive to imipenem | 0
sensitive to meropenem | 0
ascites fluid with red and white blood cells | 0
absence of pathogens in ascites fluid | 0
diagnosis of toxic epidermal necrolysis | 0
severe kidney disease | 0
vascular decompensated cirrhosis | 0
complicated diabetes mellitus type II | 0
suspected drug reaction syndrome due to carbamazepine | 0
initiation of pulse-therapy with corticosteroid | 0
topical corticosteroids | 0
topical antiseptics | 0
topical antibiotics | 0
hydro-electrolyte rebalancing | 0
continuation of basic medication | 0
favorable progress of skin lesions | 24
lack of new lesion appearance | 24
tendency of existing lesions to heal | 24
worsening of blood sugar values (499 mg/dl) | 24
worsening nitrogenous retention | 24
low alkaline reserve | 24
hyponatremia | 24
hypokalemia | 24
episode of upper gastrointestinal hemorrhage | 24
transfer to ICU | 24
satisfactory resolution of muco-cutaneous aspects | 72
reduction in corticosteroids | 72
complete discontinuation of systemic corticosteroid | 240
normalization of blood glucose levels | 240
resumption of dialysis | 240
normalization of renal function | 240
normalization of acid-base balance | 240
discharged | 360
advice to stop carbamazepine | 360
advice to stop medically related drugs | 360
