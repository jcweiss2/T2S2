19 years old | 0
male | 0
Han nationality | 0
student | 0
unmarried | 0
admitted to the hospital | 0
chest pain | -240
oliguria | -240
phlegm | -168
Nuss surgery | -6720
metal bar removal | -72
nausea | -240
vomiting | -240
repeated violent vomiting | -240
chest pain | -240
electrocardiogram | -228
ST-segment elevation | -228
coronary angiogram | -228
acute myocardial infarction | -228
myocarditis | -228
admitted to the cardiology department | -228
improved chest pain | -216
nausea | -216
vomiting | -216
anuria | -216
acute liver and renal failure | -216
transferred to the ICU | -216
emergency blood tests | -216
increased WBC | -216
neutrophiles granulocyte | -216
glutamic-pyruvic transaminase | -216
glutamic oxalacetic transaminase | -216
total bilirubin | -216
creatinine | -216
urea nitrogen | -216
serum potassium | -216
creatine kinase | -216
lactate dehydrogenase | -216
procalcitonin | -216
C-reactive protein | -216
anti-infection treatment | -216
CRRT | -216
vital signs stabilized | -216
abundant sputum | 0
difficulty in sputum expectoration | 0
CT scan | 0
left pleural effusion | 0
pericardial effusion | 0
echocardiography | 0
palpitation | 48
dyspnea | 48
sweating | 48
cyanosis | 48
heart rate | 48
blood pressure | 48
oxygen saturation | 48
intubation | 48
mechanical ventilation | 48
emergency bedside echocardiography | 48
restricted ventricular diastole | 48
stroke volume | 48
diastolic pericardial fluid | 48
thorax puncture | 48
pericardiocentesis | 48
bloody fluid | 48
coagulation function disorder | 48
coagulation factors | 48
stable | 72
fraction of inspired oxygen | 72
toxicology tests | 72
etiology tests | 72
oxygen saturation declined | 96
echocardiography | 96
pericardial effusion | 96
cardiologist | 96
thoracic surgeon | 96
radiologist | 96
chest CT | 96
sharp osteophyte | 96
Nuss surgery | 96
thoracotomy | 120
atelectasis | 120
thoracic hydrothorax | 120
pericardium | 120
pericardiotomy | 120
blood fluid | 120
scar formation | 120
horizontal mattress suture | 120
osteophytes | 120
costal osteophyte | 120
surgery | 120
drainage tube | 120
bloody fluid | 120
hemoglobin | 120
emergency surgical exploration | 120
diffuse extravasation | 120
extensive hemostasis | 120
coagulation factors | 120
mechanical ventilation | 120
anti-infection | 120
CRRT | 120
tracheotomy | 312
blood supplementing | 312
ventilator parameters | 312
antibiotics | 312
renal function recovered | 408
CRRT stopped | 408
rehabilitation exercise | 408
ventilator removed | 600
tracheal tube removed | 600
discharged | 744
follow-up | 744
normal life | 744