33 years old | 0
male | 0
admitted to the emergency department | 0
diarrhea | -24
fever | -24
vomiting stomach contents | -24
belching | -168
bloating | -168
diarrhea (past) | -168
hiatal hernia | 0
chronic nonatrophic gastritis with erosions | 0
multiple polyps in the fundus | 0
gastric polyps (0.2-0.3 cm) | 0
Yamada type II polyps | 0
fundic gland polyps | 0
colonoscopy with no abnormal findings | 0
PEG bowel preparation | -24
gastrointestinal endoscopy | 0
gastroscopy | 0
colonoscopy | 0
elevated body temperature (39°C) | 0
blood pressure 114/65 mmHg | 0
heart rate 115 beats per min | 0
respiratory rate 18 breaths per min | 0
plasma D-dimer 21800.00 μg/L | 0
BNP 7330.00 pg/mL | 0
white blood cells 35.07 × 109/L | 0
C-reactive protein 142.55 mg/dL | 0
procalcitonin 78.43 ng/mL | 0
lactic acid 3.3 mmol/L | 0
creatinine 391 μmol/L | 0
alanine aminotransferase 255 U/L | 0
aspartate aminotransferase 204 U/L | 0
total bile 72.3 μmol/L | 0
direct bile 41.1 μmol/L | 0
γ-glutamyltransferase 219 U/L |C0
abdominal CT no abnormalities | 0
lung CT small amount of inflammation in lower left lobe | 0
progressively elevated body temperature | 0
high leukocyte index | 0
metabolic acidosis | 0
respiratory rate increased to 25 breaths per min | 0
heart rate 124 beats per min | 0
blood pressure 89/60 mmHg | 0
clear systemic inflammatory response | 0
septic shock | 0
acute renal insufficiency | 0
hepatic insufficiency | 0
multiple organ failure | 0
admitted to ICU | 0
highest body temperature 40.1°C | 24
lactate level 1.0 | 48
white blood cell count 11.54 × 109/L | 48
discharged | 96
severe infection | 0
septic shock (final diagnosis) | 0
multiple organ failure (final diagnosis) | 0
good condition at 6 months postoperatively | 4320
γ-glutamyltransferase 219 U/L | 0
