36 years old | 0
male | 0
chronic smoker | 0
alcoholic | 0
admitted to the emergency ward | 0
blunt abdominal trauma | 0
resuscitation | 0
fluids | 0
norepinephrine infusion | 0
exploratory laparotomy | 0
postoperatively | 0
no oral feeds | 0
no nasogastric tube feeds | 0
central venous access | 0
parenteral nutritional support | 0
no apparent external neck swelling | 0
no neurological deficit | 0
deranged coagulation study | 0
international normalized ratio 1.8 | 0
right IJV cannulation | 0
aspirated blood | 0
aspirated white purulent color material | 0
abandoned IJV cannulation | 0
right subclavian vein cannulation | 0
cough | 2
stridor | 2
breathlessness | 2
intubated | 2
succinylcholine | 2
chest X-ray | 2
no pneumothorax | 2
transferred to Intensive Care Unit | 2
mechanical ventilation | 2
right sided subclavian CVC | 4
material aspirated | 0
detection of acid-fast bacilli | 4
Mycobacterium tuberculosis | 24
erythrocyte sedimentation rate 60 mm | 24
human immune deficiency virus positive | 24
CD4 count 180/μl | 24
X-ray chest | 24
miliary tuberculosis | 24
computed tomography of the neck | 48
retropharyngeal abscess | 48
destruction of vertebral bodies | 48
cervical brace | 48
orthopedic consultation | 48
medicine consultation | 48
pulmonary consultation | 48
category I anti-tubercular therapy | 48
cotrimoxazole tablets | 48
Pneumocystis carinii prophylaxis | 48
antiretroviral drugs | 72
tracheostomy | 168
airway compromise | -72
low-grade fever | -72
weight loss | -72
malaise | -72
night sweat | -72
vague neck pain | -72
noisy breathing | -72
respiratory distress | -72
tubercular spondylitis | -672
chronic retropharyngeal abscess | -672 
cold abscess | -672 
vertebral body destruction | -672 
abscess formation | -672 
airway spasm | 2
vagus nerve mediated laryngospasm | 2 
discharge | 720