26 years old | 0
male | 0
morbidly obese | 0
BMI 55 kg/m2 | 0
admitted to the hospital | 0
fever | -72
right lower limb pain | -72
swelling | -72
gross swelling of the entire right lower limb | 0
heart rate 111 beat per minutes | 0
temperature 38 °C | 0
leukocytosis | 0
hyperglycemia | 0
newly diagnosed with type 2 diabetes mellitus | 0
source of the infection not adequately removed | 0
extensive wound debridement | 0
above knee amputation | 72
required the use of a vasopressor | 72
acute renal failure | 0
metabolic acidosis | 0
swab culture obtained | 0
Pseudomonas aeruginosa | 0
sensitive to amikacin | 0
sensitive to gentamicin | 0
sensitive to ciprofloxacin | 0
sensitive to imipenem | 0
sensitive to meropenem | 0
sensitive to piperacillin-tazobactam | 0
sensitive to cefepime | 0
imipenem-cilastatin 500 mg every 6 h | 0
clindamycin 900 mg every 8 h | 0
daily hemodialysis | 72
septic shock | 96
multi-organ failure | 96
deteriorated | 96
death | 120
necrotizing fasciitis | 0 
tachycardia | 0
abnormal creatinine values | 0 
community-acquired P. aeruginosa | 0 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
monomicrobial necrotizing fasciitis | 0 
P. aeruginosa necrotizing infection | 0 
sub-optimal dosing of antibiotic | 0 
aggressive nature of the necrotizing infection | 0 
community-acquired | -72 
diabetes mellitus | 0 
obese patient | 0 
antibiotic dosage | 0 
treatment failure | 0 
resistance | 0 
death | 120 
acute renal failure with metabolic acidosis | 0 
sepsis | 96 
multiorgan failure | 96 
infection | -72 
necrotizing soft-tissue infection | 0 
immunocompromised patients | 0 
immunocompromised | 0 
infection sites | 0 
effectiveness of treatment | 0 
survival | 0 
diagnosis of necrotizing fasciitis | 0 
aggressive resuscitation | 0 
hemodynamic parameters | 0 
source control | 0 
surgical debridement | 0 
antimicrobial therapy | 0 
intensive patient monitoring | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
necrotizing fasciitis | 0 
infection | -72 
diabetes mellitus | 0 
obese | 0 
antibiotic | 0 
dosage | 0 
treatment | 0 
mortality | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis | 0 
P. aeruginosa infection | 0 
community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
sepsis | 96 
multiorgan failure | 96 
death | 120 
necrotizing fasciitis | 0 
infection | -72 
P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
community-acquired | -72 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 0 
infection | -72 
necrotizing fasciitis | 0 
sepsis | 96 
multiorgan failure | 96 
death | 120 
infection with community-acquired P. aeruginosa | 0 
necrotizing fasciitis caused by P. aeruginosa | 0 
P. aeruginosa | 