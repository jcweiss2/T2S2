72 years old | 0
female | 0
nonalcoholic steatohepatitis | 0
duodenal varices | 0
portosystemic encephalopathy | 0
incomplete retrograde obliteration | -1440
grade II encephalopathy | -1440
plasma ammonia level 147 µg/dL | -1440
retention rate of indocyanine green at 15 minutes 41% | -1440
hepatitis B surface antigen negative | -1440
hepatitis C virus antibody negative | -1440
antinuclear antibody negative | -1440
antimitochondrial antibody negative | -1440
huge tortuous duodenal varices | -1440
duodenal varices supplied by right colic vein | -1440
duodenal varices supplied by pancreatoduodenal vein | -1440
duodenal varices drained into inferior vena cava via right ovarian vein | -1440
spleen volume 189 mL | -1440
liver volume 595 mL | -1440
spleen/liver volume ratio 0.32 | -1440
diameter of portal vein 7.0 mm | -1440
diameter of splenic vein 6.0 mm | -1440
cobra-shaped long sheath inserted into inferior vena cava | -1440
occlusive balloon catheter inserted into right ovarian vein | -1440
obliteration of duodenal varices attempted | -1440
microcoils used | -1440
50% glucose used | -1440
absolute ethanol used | -1440
5% ethanolamine oleate with iopamidol used | -1440
incomplete obliteration of duodenal varices | -1440
encephalopathy improved to grade 0 | -1440
plasma ammonia level reduced to 39 µg/dL | -1440
febrile | -1440
drowsy | -1440
urinary incontinence | -1440
emergency admission | 0
diagnosis of recurrence of hepatic encephalopathy | 0
body temperature 39.7°C | 0
disoriented | 0
neck rigidity not evident | 0
Kernig's sign negative | 0
hemoglobin 9.7 g/dL | 0
total leukocyte count 14500/µL | 0
total platelet count 13.1 × 104/µL | 0
total bilirubin 1.3 mg/dL | 0
albumin 3.5 g/dL | 0
aspartate transaminase 37 U/L | 0
alanine transaminase 28 U/L | 0
prothrombin time 91.6% | 0
C-reactive protein 16.4 mg/dL | 0
procalcitonin 30.8 ng/mL | 0
serum ammonia 34 µg/dL | 0
Child-Pugh score 9 | 0
Child-Pugh class B | 0
mild ascites | 0
cerebral CT normal | 0
endoscopy revealed markedly reduced duodenal varices | 0
previously embolized coil partially migrated into duodenal lumen | 0
lumbar puncture | 0
purulent cerebrospinal fluid | 0
cerebrospinal fluid examination | 0
cell count 1542 /µL | 0
sugar 31 mg/dL | 0
proteins 540 mg/dL | 0
bacterial meningitis diagnosed | 0
intravenous antibiotics meropenem hydrate | 0
culture and sensitivity test of antibiotics | 120
cerebrospinal fluid culture positive for klebsiella aerogenes | 120
blood culture positive for klebsiella aerogenes | 120
urine culture positive for klebsiella aerogenes | 120
sputum culture positive for klebsiella aerogenes | 120
antibiotics changed to cefepim | 120
cefepim administered for 14 days | 120
repeat blood and cerebrospinal fluid cultures positive | 120
subsequent tests results negative | 168
trans-ileocolic vein obliteration of duodenal varices | 120
right pararectal mini-laparotomy | 120
superior mesenteric vein accessed via ileocolic vein | 120
balloon catheter inserted into right colic vein | 120
duodenal varices completely obliterated | 120
microcoils used | 120
50% glucose used | 120
portal venous pressure increased | 120
ascites increased | 120
partial splenic embolization | 288
60% infarction | 288
wedged hepatic venous pressure 23.0 cmH2O | 288
3D-CT after trans-ileocolic vein obliteration and partial splenic embolization | 360
completed embolization of duodenal varices | 360
spleen volume decreased to 85 mL | 360
liver volume increased to 889 mL | 360
corrected spleen/liver volume ratio 0.10 | 360
diameter of portal vein increased to 9.0 mm | 360
diameter of splenic vein decreased to 5.0 mm | 360
body temperature rose to 39.2°C | 600
blood culture positive for klebsiella aerogenes | 600
cefepim re-administered for 14 days | 600
blood cultures negative for bacteria | 816
neurological status regained | 816
ICG15 improved to 19% | 1008
discharged | 1008