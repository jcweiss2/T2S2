Here is the table of events and timestamps:

65 years old | 0
female | 0
history of stage IIIA lung cancer | 0
history of smoking | 0
hypertension | 0
hypothyroidism | 0
dyslipidemia | 0
spiculated suprahilar 4.5 × 2.6 cm right upper lobe (RUL) nodule | -27
multiple sub-centimeter left lung nodules | -27
lung-RADS 4X | -27
positron emission tomography/CT (PET/CT) scan | -27
adenocarcinoma | -27
stage IIIA lung adenocarcinoma | -27
T4N0M0 | -27
program death ligand-1 expression was 15% | -27
surgical resection of the mass | -27
carboplatin and paclitaxel | -27
radiation therapy | -27
repeat CT scan revealed a decrease in the RUL mass | -12
adjuvant immunotherapy with durvalumab | -12
pneumonitis | -12
staging chest CT showed an increase in the RUL mass | -6
further follow-up chest CT showed an increase in the RUL mass | -6
routine follow-up by the pulmonary medicine clinic | -6
abdominal and pelvic CT scan | -6
no distant metastasis | -6
stable lung nodules | -6
5 subsequent chest CT scans | -6
last chest CT scan in June 2022 | -6
abdominal pain | -6
pancreatic head lesion | -6
PET/CT scan | -6
fluorodeoxyglucose-avid mass in the pancreatic head | -6
SUV max of 13.3 | -6
increased uptake in the porta hepatis | -6
no other regions of metastases | -6
no lymphadenopathy | -6
brain MRI scan | -6
negative for intracranial metastasis | -6
palliative radiation therapy to the pancreatic mass | -6
combination chemotherapy with carboplatin and pemetrexed | -6
3 cycles completed | -6
electrolyte derangements | -6
acute anemia | -6
hemoglobin nadir of 6.9 g/dL | -6
transfusion | -6
new 9 mm left lower lobe nodule | -6
staging PET/CT scan | -6
decreased metabolic activity in the pancreatic mass | -6
metabolic activity in the new left lower lobe nodule | -6
uncertainty regarding treatment continuation | -6
no further treatments | -6
rapid response called | -3
saturating at 87% on 3 L of oxygen via nasal cannula | -3
using her accessory muscles | -3
blood pressure of 84/70 | -3
heart rate of 138 | -3
increased dyspnea | -3
cough | -3
generalized weakness | -3
imaging studies on admission | -3
right lung consolidation concerning for an infectious process | -3
loculated pleural effusion | -3
treatment for acute hypoxic respiratory failure in the context of sepsis secondary to pneumonia | -3
broad-spectrum antibiotics | -3
oxygen supplementation | -3
bilevel-positive airway pressure | -3
episode of altered mentation and worsening hypoxemia | -3
critical care consult | -3
vasopressor support | -3
palliative medicine team consulted | -3
transition to inpatient hospice care | -3
inpatient hospice care | -3
passed peacefully under comfort measures | -3