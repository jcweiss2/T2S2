80 years old | 0
female | 0
Alzheimer’s dementia | 0
diabetes mellitus | 0
hypertension | 0
chronic kidney disease | 0
admitted to the ICU | 0
hypotension | 0
lactic acidosis | 0
progressive altered mental status | -336
physical decline | -336
initial blood pressure 89/56 | 0
normal heart rate | 0
oxygen saturation normal | 0
no fever | 0
no tachypnea | 0
lactic acid 3.6 mmol/L | 0
leukocytosis | 0
neutrophilic predominance | 0
troponin peaked at 1104 pg/mL | 0
Wells score 0 points | 0
D-dimer not obtained | 0
treated with fluids | 0
treated with broad-spectrum antibiotics | 0
blood pressure improved | 24
lactic acidosis resolved | 24
troponin elevation secondary to demand ischemia | 24
blood cultures negative | 24
transferred to the gerontology unit | 48
afebrile | 48
heart rate 80 | 48
blood pressure 117/62 | 48
SpO2 99% on room air | 48
jugular venous distension | 48
normal cardiopulmonary auscultatory exam | 48
no peripheral edema | 48
no asymmetric lower extremity swelling | 48
dilated RV with akinesis of the mid-RV free wall | 48
McConnell’s sign | 48
diastolic septal flattening | 48
D-sign | 48
dilated IVC with minimal inspiratory variation | 48
S1Q3T3 pattern on ECG | 48
D-dimer 51,190 ng/mL | 48
saddle PE involving both main pulmonary arteries | 48
RV strain on CT angiography | 48
initiated on heparin infusion | 48
transitioned to oral apixaban | 72
taking megestrol as an outpatient | -720
discharged | 168