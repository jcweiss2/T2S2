85 years old | 0
female | 0
admitted to the hospital | 0
chest pain | -72
dyspnea | 0
hypertension | -672
dyslipidemia | -672
elevated troponin T level | 0
ST depression in V2–5 | 0
pulmonary congestion | 0
severe mitral regurgitation | 0
P2 prolapse | 0
99% stenosis of the mid-portion of the left circumflex artery | 0
intra-aortic balloon pumping | 0
intubated | 0
transesophageal echocardiography | 0
papillary muscle rupture | 0
cardiogenic shock | 0
inotrope support | 0
emergency PCI | 12
MICS-MVR | 12
cardiopulmonary bypass | 12
cardiac arrest | 12
antegrade cardioplegia | 12
mitral valve replacement | 12
discontinued intra-aortic balloon pumping | 24
extubated | 48
sepsis | 96
antibacterial treatment | 96
discharged from the ICU | 144
postoperative TTE | 144
normal cardiac and bioprosthetic valve function | 144
walk 200 m independently | 144
transferred to another hospital | 144