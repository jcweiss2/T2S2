72 years old | 0
male | 0
mechanical fall | -72
lying on the floor for 3 days | -72
Stage IVA (T2N2bM0) squamous cell carcinoma (positive HPV) of bottom of tongue | -5760
completed concurrent chemoradiotherapy with cetuximib and radiotherapy | -5760
weakness | 0
pain in right wrist | 0
pain in left hip | 0
epiphora | 0
pain in left eye | 0
limited range of motion of both hips | 0
minimal erythema | 0
palpable trace effusion | 0
tenderness to palpation over dorsal distal radius | 0
tenderness to palpation over volar wrist | 0
tenderness to palpation over carpus on right hand and wrist | 0
left eye matted eyelashes | 0
mucopurulent conjunctival secretions | 0
corneal edema | 0
hypopyon with fibrinous membrane in pupil | 0
no red glow seen | 0
pupil fixed and non-reactive | 0
white blood cell count of 6.6 K/cmm | 0
thrombocytopenia (platelet count of 47.0 K/cmm) | 0
renal impairment (blood urea nitrogen of 47.0 mg/dL; creatinine of 1.4 mg/dL) | 0
procalcitonin 5.13 ng/mL | 0
blood cultures growth of Gram-positive cocci in chains | 0
beta-hemolytic Group C Streptococcus dysgalactiae subsp. equisimilis identified | 0
left eye pain | 0
left eye watering | 0
decreased vision in left eye | 0
B scan ultrasound of the left eye showed vitreous debris | 0
aqueous tap of left eye | 0
vitreous tap of left eye | 0
intravitreal injection of vancomycin and ceftazidime | 0
vitreous culture growth of Gram-positive Streptococcus dysgalactiae subsp. equisimilis | 0
transthoracic echocardiography (TTE) at day 3 showed bicuspid aortic valve with mild to moderate aortic regurgitation | 72
TTE at day 3 showed normal left ventricular function | 72
TTE at day 3 showed mild to moderate dilatation | 72
TTE at day 3 showed normal right ventricular size and function | 72
TTE repeat at day 6 showed aortic valve vegetation | 144
TTE repeat at day 6 could not exclude abscess or anterior mitral valve leaflet vegetation | 144
transesophageal echocardiography (TEE) at day 9 showed small, mobile vegetation on the non-coronary cusp of the aortic valve | 216
TEE at day 9 showed thickened aortic root | 216
TEE at day 9 showed echodensity in the posterior aspect of the aortic root adjacent to the right atrium | 216
TEE at day 9 showed moderate aortic valve vegetation | 216
TEE at day 9 noted thickened mitral valve suggesting possible microperforation | 216
TEE at day 9 showed mobile echodensity on the posterior mitral valve (0.3 × 0.5 cm) | 216
TEE at day 9 showed mild-moderate mitral valve regurgitation | 216
treated with intravenous vancomycin every 12 hours for 2 days | 0
followed by intravenous penicillin G every 4 hours | 48
diagnosed with infective endocarditis (IE) using modified Duke criteria | 0
left eye vision worsened to light perception | 0
received another intravitreal injection in left eye | 0
treated with topical trimethoprim/sulfamethoxazole | 0
treated with topical prednisolone acetate | 0
treated with topical atropine | 0
scheduled for vitrectomy of left eye | 0
no light perception in left eye | 0
vitrectomy cancelled | 0
orthopedic service ruled out septic arthritis | 0
right humerus showed no evidence of fracture or dislocation | 0
right wrist showed no evidence of fracture or dislocation | 0
right hand showed no evidence of fracture or dislocation | 0
right shoulder showed no evidence of fracture or dislocation | 0
no soft tissue swelling | 0
magnetic resonance imaging of thoracic and lumbar spine with contrast showed no evidence of infection | 0
otolaryngologists found no infection or new lesions on ear, nose, and throat | 0
all blood cultures negative during treatment | 0
transferred to another facility for aortic valve replacement | 0
acute heart failure secondary to worsening aortic regurgitation | 0
developed hypoxic respiratory distress | 0
chest x-ray showed pulmonary edema | 0
temporarily placed on BiPAP | 0
started on dobutamine | 0
bicuspid aortic valve replaced with prosthetic valve | 24
aortic root abscess debrided | 24
transferred to general medicine floor after 3 days | 72
died | unknown
underwent valve replacement | 24
loss of vision | 0
myocardial abscess | 216
endophtalmitis | 0
infective endocarditis | 0
