19 years old | 0
male | 0
army officer | 0
admitted to the hospital | 0
fever | -120
arthralgia | -120
myalgia | -120
headache | -120
productive cough | -120
yellowish sputum | -120
chest heaviness | -120
dyspnea | -120
diarrhea | -120
reduced oral intake | -120
no history of travelling | 0
no recent jungle activities | 0
no past medical illness | 0
no previous hospitalization | 0
no medical treatment for current condition | 0
conscious | 0
dehydrated | 0
cold peripheries | 0
febrile | 0
temperature of 38.5°C | 0
hypotensive | 0
blood pressure of 81/53 mmHg | 0
tachycardic | 0
146 beats per minute | 0
tachypnoeic | 0
30 breaths per minute | 0
oxygen saturation of 75-80% | 0
coarse crepitation over both lower zone of lungs | 0
tenderness at epigastric region | 0
palpable liver | 0
no cervical lymph nodes | 0
no inguinal lymph nodes | 0
no axillary lymph nodes | 0
haemoglobin of 11.3 g/dL | 0
low white blood cell count | 0
neutrophil predominance | 0
platelet count of 80 × 10^6/L | 0
C-reactive protein of 28.28 mg/dL | 0
acute kidney injury | 0
serum sodium of 137 mmol/L | 0
serum potassium of 3.7 mmol/L | 0
serum urea of 14 mmol/L | 0
serum creatinine of 206 μmol/L | 0
liver function tests normal | 0
serum albumin of 22 g/dL | 0
creatinine kinase of 351 IU/L | 0
arterial blood gases on room air | 0
pH of 7.378 | 0
pCO2 of 37 mmHg | 0
pO2 of 52.7 mmHg | 0
O2 saturation of 89% | 0
HCO3 of 21.7 mmol/L | 0
Dengue NS-1 Antigen negative | 0
IgG and IgM antibody negative | 0
chest radiograph showed consolidation | 0
diagnosis of severe community acquired pneumonia | 0
acute kidney injury | 0
resuscitated with normal saline | 0
started on non-invasive ventilation | 0
inotropic support | 0
commenced empirically with ceftriaxone and azithromycin | 0
intubation and mechanical ventilation | 24
bronchoscopy on day 2 | 48
copious amount of haemoserous and greenish secretion | 48
repeated chest radiograph showed worsening consolidation | 48
antibiotics upgraded to meropenem and cloxacillin | 48
antiviral oseltamivir added | 48
continuous venous-venous haemofiltration | 48
severe metabolic acidosis | 48
oliguric acute kidney injury | 48
persistent spiking of temperature | 48
worsening of septic parameters | 48
refractory hypotension | 48
maximum dose of multiple inotropic agents | 48
patient succumbed | 72
blood cultures negative | 72
atypical bacterial and Leptospiral serologies negative | 72
Hepatitis B/C and HIV serologies undetected | 72
respiratory viruses screening negative | 72
tracheal aspiration and bronchoalveolar lavage positive for MDR Acinetobacter baumannii | 72
MDR Acinetobacter baumannii susceptible only to polymyxin B | 72
minimum inhibitory concentration of 0.5 μg/ml | 72
MDR Acinetobacter baumannii resistant to penicillin group | 72
ampicillin/sulbactam | 72
third generation cephalosporins | 72
fluoroquinolone | 72
carbapenem group | 72
PCR for carbapenemases genes NDM, OXA-23, OXA 24 or OXA-58 not performed | 72