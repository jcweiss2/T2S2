56 years old | 0
male | 0
admitted to the hospital | 0
infection around the limbs of an aortic bifurcation graft | 0
large abscess in the right groin | 0
severe systemic inflammatory response | 0
physiologic severe systemic inflammatory response | 0
biochemical severe systemic inflammatory response | 0
aortobifemoral graft | -2400
lifestyle-limiting claudication | -2400
exercise tolerance of 50 yards | -2400
medication controlled hypertension | -2400
previous transient ischemic attack | -3600
acute occlusion of the left limb of the graft | -1200
thrombectomize the limb of the aortic bifurcation graft | -1200
femoral crossover graft | -1200
clinical outcome from this treatment was good | -1200
acute right groin pain | -600
swelling | -600
erythema | -600
abscess identified on a computed tomography (CT) scan | -600
Proteus mirabilis | -600
Staphylococcus epidermidis | -600
Enterococcus faecalis | -600
intravenous daptomycin | -600
teicoplanin | -600
oral ciprofloxacin | -600
surgical re-exploration | -600
inflammatory fluid and tissue identified at the aortic anastomosis | -600
explant of the aortobifemoral graft | -600
explant of the femoral crossover graft | -600
rifampicin-bonded graft | -600
omental wrap | -600
severe systemic inflammatory response with pyrexia | 0
tachycardia | 0
large right groin abscess | 0
anterior abdominal wall and groin cellulitis | 0
CT angiography | 0
large collection in the right groin | 0
inflammatory changes seen to the level of the aortic anastomosis | 0
inflammatory changes seen around the left limb of the graft | 0
patent native right common iliac artery | 0
patent distal aorta | 0
patent common femoral arteries | 0
patent profunda femoris arteries | 0
occluded right superficial femoral artery | 0
severe stenosis at the adductor hiatus | 0
surgical options considered | 0
decision made to proceed with NAIS | 0
small bowel fistulae onto the graft | 0
duodenum to the main body of the graft | 0
distal ileum to the right limb of the graft | 0
infrarenal aortic clamp | 0
Dacron graft completely excised | 0
arteriosclerosis of the aortic wall | 0
aortic anastomosis | 0
previous aortotomy | 0
distal anastomoses to the common femoral arteries | 0
sartorius flaps performed on both sides | 0
vasopressor support | 24
renal replacement therapy | 24
organ dysfunction | 24
sepsis | 24
major surgery | 24
lower limb ischemia/reperfusion injury | 24
four-compartment fasciotomy of the left leg | 48
compartment syndrome | 48
ischemia/reperfusion | 48
venous hypertension | 48
deep venous harvest | 48
severe abdominal pain | 264
back pain | 264
hypovolemic shock | 264
CT angiogram | 264
large, contained false aneurysm at the aortic anastomosis | 264
endovascular salvage | 264
left axillary artery surgically exposed | 264
directly punctured | 264
GORE Dry Seal sheath | 264
stiff wire | 264
suprarenal aorta | 264
Amplatzer vascular plugs | 264
native right common iliac artery occluded | 264
distal aorta occluded | 264
Medtronic flared limb | 264
caliber mismatch | 264
native aorta | 264
deep vein | 264
flared stent graft | 264
completion angiography | 264
exclusion of the pseudoaneurysm | 264
discharged | 360
intravenous ertapenem | 360
daptomycin | 360
multidrug-resistant E coli | 360
vancomycin-resistant Enterococcus | 360
oral doxycycline | 360
trimethoprim | 360
white cell count | 2160
C-reactive protein | 2160
albumin | 2160
surveillance CT angiogram | 2160
inflammatory change around the aortic reconstruction | 2160