39 years old | 0
male | 0
admitted to the hospital | 0
skin flare-up | -168
tenderness in the right upper limb | -168
scratches on the right upper arm | -168
minor abrasion | -168
sore throat | -96
fever | -96
erythema | 0
swelling of the right upper arm | 0
swelling of the right lateral thorax | 0
pain | 0
no paralysis | 0
no contracture of the right hand or wrist | 0
increased white blood cell count | 0
increased neutrophils | 0
decreased hemoglobin | 0
decreased platelet | 0
elevated C-reactive protein | 0
decreased total protein | 0
decreased albumin | 0
elevated aspartate aminotransferase | 0
elevated alanine aminotransferase | 0
elevated total bilirubin | 0
elevated creatine kinase | 0
elevated blood urea nitrogen | 0
elevated creatinine | 0
decreased sodium | 0
decreased potassium | 0
decreased chloride | 0
normal glucose | 0
elevated presepsin | 0
elevated prothrombin time | 0
elevated fibrinogen | 0
decreased antithrombin 3 | 0
computed tomography findings | 0
LRINEC score of 9 | 0
shock | 0
tachypneic state | 0
noradrenaline infusion | 0
vasopressin infusion | 0
administration of meropenem | 0
administration of vancomycin | 0
administration of clindamycin | 0
tracheal intubation | 0
ventilatory assistance | 0
emergency surgery | 0
incision in the dorsal triceps brachii | 0
excision of the fascia | 0
contamination of latissimus dorsi and triceps brachii | 0
presence of pus | 0
no contamination of the right forearm | 0
transfer to intensive care unit | 0
positive blood cultures for Streptococcus pyogenes | 0
positive drainage cultures for Streptococcus pyogenes | 0
flare of the right precordia exacerbated | 96
incision from precordia to medial elbow | 96
debridement of contaminated tissues | 96
marking nerves and vessels with vessel tapes | 96
open wounds | 96
daily wound cleaning | 96
fasciotomy on hospitalization days 5 and 6 | 120
transfer to ward | 168
administration of ampicillin | 216
administration of clindamycin | 216
daily wound cleaning in ward | 216
detection of Klebsiella aerogenes | 360
change to cefepime | 360
thorough debridement on day 19 | 456
identification of nerves and vessels | 456
wound closure with skin graft | 1080
discharge | 1944
administration of cefepime until day 36 | 864
administration of oral minocycline | 1944
no nerve injuries at 12 months | 8760
active shoulder ROM | 8760
active elbow ROM | 8760
active forearm ROM | 8760
no ROM limitations in wrist and fingers | 8760
hypertrophic scar contracture | 8760
