75 years old | 0  
    male | 0  
    hypertension | 0  
    sequelae of ischemic stroke | 0  
    mild right hemiplegia | 0  
    fell into a creek | -144  
    face submerged in water | -144  
    rescued | -144  
    brought to local hospital | -144  
    Glasgow Coma Scale E3V3M6 | -144  
    body temperature 33.4°C | -144  
    heart rate 88 beats/min | -144  
    blood pressure 120/60 mmHg | -144  
    respiratory rate 26 breaths/min | -144  
    oxygen saturation 92% | -144  
    no obvious injury | -144  
    bilateral coarse crackles | -144  
    hypothermia | -144  
    rewarming using warming blanket | -144  
    antibiotic therapy (ampicillin and sulbactam) | -144  
    non-invasive ventilation | -144  
    oxygenation deteriorated to 80% | -144  
    intubated | -144  
    mechanically ventilated | -144  
    transferred to tertiary hospital | -144  
    sedated with propofol | 0  
    body temperature 36.4°C | 0  
    heart rate 104 beats/min | 0  
    blood pressure 123/84 mmHg | 0  
    respiratory rate 30 breaths/min | 0  
    oxygen saturation 91% | 0  
    bilaterally diminished breath sounds | 0  
    arterial blood gas pH 7.34 | 0  
    PaCO2 42 mmHg | 0  
    PaO2 199 mmHg | 0  
    HCO3 21.9 mmol/L | 0  
    white blood cell count 2980/μL | 0  
    neutrophils 63.5% | 0  
    hemoglobin 15.3 g/dL | 0  
    platelet 159,000/μL | 0  
    C-reactive protein 0.6 mg/dL | 0  
    procalcitonin 59.37 ng/mL | 0  
    normal ejection fraction | 0  
    no valvular disease | 0  
    chest radiography diffuse infiltrates | 0  
    CT diffuse infiltrates | 0  
    no pleural effusion | 0  
    diagnosis of ARDS | 0  
    aspiration pneumonitis | 0  
    septic shock | 0  
    treated with isotonic crystalloids | 0  
    meropenem 1.0 g every 12 hrs | 0  
    vasopressors | 0  
    protective ventilation | 0  
    methylprednisolone 80 mg daily started | 72  
    beta-D-glucan elevated 37.6 pg/mL | 96  
    vasopressors stopped | 120  
    hypoxia did not improve | 120  
    tracheal aspirate culture positive Aeromonas hydrophila | 144  
    blood culture negative | 144  
    switched to piperacillin/tazobactam | 144  
    hypoxia worsened | 168  
    died | 168  
    autopsy CT diffuse infiltrates | 168  
    lungs congested | 168  
    pulmonary embolus right pulmonary artery | 168  
    no femoral vein embolus | 168  
    Grocott staining diffuse filamentous fungi | 168  
    fungi identified Aspergillus fumigatus | 168  
    invasive aspergillosis | 168  
    pulmonary embolism | 168  
    fungi in heart | 168  
    fungi in stomach | 168  
    fungi in thyroid gland | 168  
    no focal brain lesion | 168  
    no history of aspiration pneumonia | 0  
    good swallowing function | 0  
    no co-morbidities except hypertension | 0  
    elevated β-glucan misinterpreted | 96  
    no galactomannan measurement | 0  
    primary hospital culture positive Aspergillus fumigatus | 168  
    no bronchoscopy performed | 0  
    no BAL performed | 0  
    long history of smoking | 0  
    impaired ciliary activity | 0  
    hypothermia at presentation | -144  
    low white cell count | 0  
    methylprednisolone use worsened aspergillosis | 72  
    thromboprophylaxis with heparin | 0  
    compression stockings | 0  
    no antifungal therapy administered | 168  
    no antifungal therapy considered | 0  
    no invasive procedures | 0  
    rapid disease progression | 168  
    severe hypoxia | 0  
    pulmonary embolism caused by angioinvasiveness | 168  
    no COPD history | 0  
    impaired immune response | 0  
    no survivors with CNS infection | 168  
    length of stay 7 days | 168  

    <|eot_id|>
    