68 years old | 0
    male | 0
    admitted to ICU | 0
    hypoxemic respiratory failure | -24
    septic shock | -24
    trachea intubated | -24
    fluid resuscitation | -24
    vasopressor support | -24
    right IJV CVC insertion | -24
    acute renal failure | -24
    anuria | -24
    metabolic acidosis (HCO3 12 mEq/L) | -24
    hyperkalemia (K+ 6.8 mEq/L) | -24
    hemodialysis planned | -24
    left IJV chosen for dialysis catheter | -24
    right IJV already catheterized | -24
    femoral vein higher risks (infection, thrombosis, occlusion) | -24
    positioning with head slightly lower | 0
    left neck cleaned with chlorhexidine | 0
    draped | 0
    Seldinger technique under ultrasound guidance | 0
    local anesthesia (4 ml 2% lignocaine) | 0
    IJV located with ultrasound | 0
    vein punctured at 45° angle | 0
    free aspiration of blood confirmed | 0
    guidewire threaded | 0
    resistance after 5 cm guidewire | 0
    guidewire removed | 0
    syringe connected for free blood aspiration | 0
    needle in vein confirmed | 0
    reattempted guidewire insertion | 0
    resistance again after 5 cm | 0
    normal breath sounds | 0
    normal respiratory rate | 0
    oxygen saturation 98% | 0
    no subcutaneous emphysema | 0
    no hematoma | 0
    no venous congestion | 0
    no limb ischemia | 0
    senior ICU registrar called | 0
    guidewire and needle scanned | 0
    guidewire inside vein | 0
    loop visualized (dual-point echogenicity) | 0
    introducer needle retracted | 0
    guidewire pulled back under ultrasound | 0
    loop disappeared | 0
    guidewire advanced caudally | 0
    dilation | 0
    dialysis catheter railroaded | 0
    guidewire removed | 0
    correct placement confirmed with USG | 0
    blood aspirated in both ports | 0
    free flow confirmed | 0
    chest X-ray performed | 24
    carcinoma of pyriform fossa | -672
    no comorbidities | -672
    hemodialysis catheter successfully placed | 24
    