42 years old | 0
female | 0
admitted to the hospital | 0
motorcycle accident | -336
fracture of the middle third of the right clavicle | -336
Allman's group I | -336
AO 15-B1 | -336
deviation >2 cm | -336
right shoulder abrasions | -336
prescribed analgesics | -336
no orientation regarding the use of a sling | -336
no need for therapeutic follow-up with a specialist | -336
pain | -336
fever | -336
local hyperemia | -336
hospitalization | -336
febrile peaks | -336
local edema | -336
skin fluctuation on the right clavicle region | -336
drainage of a purulent secretion | -336
abscess drainage | -336
cleansing with 0.9% saline solution | -336
leukogram presented a WBC of 12,000/mm3 | -336
ESR: 25 mm/h | -336
CRP: 11 mm/dl | -336
intravenous antibiotic therapy | -336
ceftriaxone 1 g 12/12 h | -336
metronidazole 500 mg 8/8 h | -336
clindamycin 600 mg 8/8 h | -336
admitted to this medical service in Salvador, Bahia State | -600
extensive lesion of the right hemithorax | -600
toxemia | -600
sepsis | -600
clavicle bone exposure | -600
extensive necrosis of the skin | -600
no neurovascular alterations | -600
leukogram presented with 21,000 WBC/mm3 | -600
ESR: 44 mm/h | -600
PCR: 20 mm/dl | -600
creatinine: 1.3 mg/dl | -600
urea: 48 mg/dl | -600
CPK: 900 u/l | -600
magnetic resonance imaging (MRI) of the thorax | -600
inflammatory process in the anterior region of the thorax | -600
admitted to the intensive care unit (ICU) | -600
infectious diseases team requested surgical debridement | -600
modified antibiotic therapy | -600
meropenem 1 g 8/8 h | -600
vancomycin 1 g 12/12 h | -600
anti-tetanus prophylaxis | -600
surgical debridement | -576
right clavicle resection | -576
aggressive debridement of the devitalized tissue | -576
soft tissue and bone cultures were collected | -576
important clinical improvement | -576
discharged from the ICU | -552
reduction of the WBC and inflammatory markers | -552
purulent secretion diminished | -552
special dressing | -528
borders of the lesion ceased to evolve with necrosis | -528
raw area was without purulent secretion | -528
forming granulation tissue | -528
final bone and soft tissue culture results were negative | -528
skin graft | -432
normal laboratory tests | -432
evolved without new signs of infection | -432
discharged from the hospital | -432
wound presented complete healing | -240
excellent upper limb functional score | -240
UCLA score: 33 points | -240
Constant Score: 93 points | -240