39 years old | 0
female | 0
ovarian cancer | -336
stage III | -336
TAH with BSO | -336
paclitaxel | -240
carboplatin | -240
melena | -192
hematochezia | -192
abdominal tenderness | -192
rebound tenderness | -192
neutropenia | -192
high fever | -192
tachypnea | -192
hypotension | -192
cyanosis | -192
neutropenic/septic shock | -192
ascending colon perforation | -192
emergent total colectomy | -192
intubated | -192
alert and oriented | -192
difficulty in weaning from mechanical ventilation | -168
severe tachypnea | -168
labored breathing | -168
midazolam | -168
G-CSF injection | -168
ANC less than 50/µl | -168
chemotherapy induced neutropenia | -168
sepsis | -168
G-CSF | -168
antibiotics | -168
Piperacillin/tazobactam | -168
midazolam stopped | -120
extubated | -120
dyspnea | -120
deteriorating levels of consciousness | -120
reintubation | -96
brain CT | -96
EEG | -96
no abnormal findings | -96
partial seizure | -48
GTC seizure | -48
seizure controlled | -48
midazolam | -48
ativan | -48
phenytoin | -48
diffuse brain swelling | -24
severe diffuse cerebral dysfunction | -24
hyperammonemia | -24
respiratory alkalosis | -24
metabolic alkalosis | -24
sodium benzoate | -24
mannitol | -24
recurrent episodes of GTC seizure | 0
status epilepticus | 0
desaturation | 24
hypotension | 24
death | 48