66 years old | 0
male | 0
dual-chamber pacemaker | -13104
sick sinus syndrome | -13104
paroxysmal atrial fibrillation | -13104
severe lumbar back pain | 0
mental status changes | 0
hypotension | 0
acute renal failure | 0
hypoxemic respiratory failure | 0
emergent intubation | 0
severe sepsis | 0
hemodynamic support | 0
vasopressin | 0
norepinephrine | 0
blood cultures | 0
methicillin-sensitive Staphylococcus aureus | 0
vancomycin | 0
nafcillin | 0
transthoracic echocardiogram | 0
left ventricular ejection fraction | 0
patent foramen ovale | 0
Doppler of the intra-atrial septum | 0
computed tomography scan | 0
osteomyelitis | 0
magnetic resonance imaging | 0
septic emboli | 0
transesophageal echocardiogram | 0
vegetation | 0
right atrium | 0
pacemaker lead | 0
tricuspid valve | 0
right ventricle | 0
cardiothoracic surgery | 0
surgical intervention | 0
laser lead extraction | 0
Indigo Thrombectomy System | 0
intracardiac echocardiography | 0
vacuum-assisted vegetation removal | 0
femoral veins | 0
GORE DrySeal Flex introducer sheath | 0
CARTO SoundStar | 0
Indigo CAT8 XTORQ | 0
aspiration | 0
vegetation extraction | 0
lead extraction | 0
pocket inspection | 0
suture | 0
hemostasis | 0
figure-of-8 closures | 0
pathology | 0
gram-positive cocci | 0
methicillin-sensitive Staphylococcus aureus | 0
tissue necrosis | 48
lactic acidosis | 48
worsening renal failure | 48
withdraw care | 72
extubation | 72
death | 72