80 years old | 0
male | 0
admitted to the hospital | 0
hypotension | 0
denied chest pain | 0
denied shortness of breath | 0
denied fever | 0
denied cough | 0
denied palpitation | 0
denied nausea | 0
denied vomiting | 0
denied abdominal pain | 0
denied changes in urinary habits | 0
denied changes in bowel habits | 0
WBC count 16.5 K/UL | 0
Hgb 14.3 GM/DL | 0
PLT 115 K | 0
Creatinine 12.59 MG/DL | 0
BUN 56 MG/DL | 0
Sodium 133 MMOL/L | 0
Potassium 5.4 MMOL/L | 0
BNP 143 PG/ML | 0
Troponin 0.05 NG/ML | 0
EKG ST segment elevation V3, V4, V5 | 0
EKG Q wave II, III, AVF | 0
diagnosed with acute STEMI | 0
aspirin 325 mg | 0
clopidogrel 300 mg | 0
atorvastatin 80 mg | 0
heparin 3500 units/kg | 0
cardiac catheterization | 0
coronary angiography chronic total right coronary artery occlusion | 0
collaterals from left | 0
left coronary arteries patent | 0
left ventriculography mid to apical akinesis | 0
left ventriculography basal hyperkinesis | 0
transferred to ICU | 0
levophed started | 0
CK-MB 11.6 ng/ml | 4
Troponin 2.10 | 4
EKG resolution ST elevation anterior leads | 6
leukocytosis | 0
septic shock | 0
cardiogenic shock | 0
vancomycin started | 6
Zosyn started | 6
transthoracic echocardiography LVEF 25-30% | 12
elevated LV end diastolic pressure | 12
akinesis left and right ventricles | 12
remained chest pain free | 12
continued levophed | 12
neosynephrine started | 12
sepsis workup unremarkable | 24
repeat echocardiogram LV thrombus | 24
akinesis both ventricles | 24
anticoagulation heparin started | 24
plan repeat echo 3-4 days | 24
hemodynamically unstable | 72
died | 72
autopsy not performed | 72
peripheral artery disease | -Infinity
hypertension | -Infinity
end stage renal disease | -Infinity
peritoneal dialysis | -Infinity
nursing home | -Infinity
