71 years old | 0
male | 0
Japanese | 0
admitted to the hospital | 0
right upper quadrant abdominal pain | -168
exacerbation of chronic diarrhea | -120
fever | -48
headache | -48
disturbance of consciousness | -48
birthplace was the Amami Islands in Japan | 0
frequently visited Okinawa in his childhood | 0
frequent travel to the Solomon Islands on business | -1440
hepatitis B virus carrier | 0
HTLV-1 carrier | 0
chronic alcohol abuse | 0
temperature of 36.0 ℃ | 0
blood pressure of 117/85 mmHg | 0
pulse rate of 95 beats per minute | 0
respiratory rate of 24 per minute | 0
oxygen saturation of 94% | 0
neck rigidity | 0
whole abdominal pain | 0
severe thrombocytopenia | 0
elevated liver enzyme levels | 0
liver abscess | 0
meropenem administration | 0
intensive care | 0
respirator support | 0
deteriorated mental status | 0
blood culture revealed K. pneumoniae | 96
cerebrospinal fluid culture revealed K. pneumoniae | 96
direct microscopy of the stool showed rhabditiform larvae of S. stercoralis | 96
ivermectin administration | 96
coma | 96
discontinuation of sedation drugs | 96
electroencephalogram revealed flat brain waves | 144
head CT revealed pseudo-subarachnoid hemorrhaging signs | 144
severe cerebral edema | 144
cardiopulmonary arrest | 168
death | 168
autopsy | 168
necrosis with neutrophil infiltration in the liver tissue | 168
neutrophil infiltration in the meninges and cerebral parenchyma | 168
rhabditiform larvae of S. stercoralis in the cecum polyp | 168
no S. stercoralis larvae in the liver or brain tissue | 168
polyp in the cecum | 168
chronic strongyloidiasis | 0
hypermucoviscous K. pneumoniae infection | 0
K1 capsular serotype | 0
ST23 sequence type | 0
positive for magA, rmpA, iutAfimH, aerobactin, and iroN | 0