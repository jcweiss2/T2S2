39 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
palpable mass on right breast | -168 | 0 | Factual
Hodgkin lymphoma | -6336 | -6336 | Factual
chemotherapy | -6336 | -6336 | Factual
mantle field radiation | -6336 | -6336 | Factual
inflammatory colitis | -6336 | -168 | Factual
mesalazine | -168 | -168 | Factual
family history of myxoid liposarcoma | 0 | 0 | Factual
no family history of breast or ovarian tumors | 0 | 0 | Factual
radiological examination of breast | -168 | 0 | Factual
invasive ductal carcinoma | -168 | 0 | Factual
triple-negative phenotype | -168 | 0 | Factual
MIB1 85% | -168 | 0 | Factual
staging CT scan | -168 | 0 | Factual
no distant metastasis | -168 | 0 | Factual
neoadjuvant chemotherapy | -168 | 0 | Factual
paclitaxel | -168 | 0 | Factual
carboplatin | -168 | 0 | Factual
first cycle of chemotherapy | -120 | -96 | Factual
no hematological toxicity | -96 | 0 | Factual
port-à-cath insertion | -96 | -96 | Factual
fever | -72 | -72 | Factual
subcutaneous cellulitis | -72 | -72 | Factual
colliquative necrosis | -72 | -72 | Factual
elevated white blood cell count | -72 | -72 | Factual
neutrophilia | -72 | -72 | Factual
elevated C-reactive protein | -72 | -72 | Factual
broad-spectrum i.v. antibiotic therapy | -72 | -72 | Factual
piperacillin/tazobactam | -72 | -72 | Factual
daptomycin | -72 | -72 | Factual
PORT rimotion | -72 | -72 | Factual
necrosectomy | -72 | -72 | Factual
defervescence | -48 | -48 | Factual
improvement in subcutaneous cellulitis | -48 | -48 | Factual
improvement in blood works | -48 | -48 | Factual
new febrile seizure | -48 | -48 | Factual
WBC rise | -48 | -48 | Factual
worsening of skin lesion | -48 | -48 | Factual
second necrosectomy | -48 | -48 | Factual
peripheral blood cultures negative | -48 | -48 | Factual
skin plug negative | -48 | -48 | Factual
i.v. catheter tip positive for Klebsiella pneumoniae | -48 | -48 | Factual
antibiotic therapy modified | -48 | -48 | Factual
chest/abdomen CT scan | -48 | -48 | Factual
mediastinitis | -48 | -48 | Factual
bilateral pleural effusion | -48 | -48 | Factual
left pulmonary atelectasis | -48 | -48 | Factual
thoracoscopy | -48 | -48 | Factual
pleural and mediastinal drainage | -48 | -48 | Factual
sepsis | -48 | 0 | Factual
broad-spectrum antibiotic and antifungal therapy | -48 | 0 | Factual
hemodynamic support | -48 | 0 | Factual
non-invasive ventilation | -48 | 0 | Factual
specimens of skin and subcutaneous and muscular tissue analyzed | -48 | -48 | Factual
intensive inflammatory infiltrate | -48 | -48 | Factual
neutrophils | -48 | -48 | Factual
differential diagnosis included PG | -48 | -48 | Factual
systemic methylprednisolone | -24 | 0 | Factual
topical cyclosporine | -24 | 0 | Factual
seriate chest X-ray and CT scan | -24 | 0 | Factual
progressive resolution of mediastinitis | -24 | 0 | Factual
progressive resolution of pleural effusion | -24 | 0 | Factual
wound improvement with scar | -24 | 0 | Factual
blood works indicated progressive normalization | -24 | 0 | Factual
breast ultrasound | 0 | 0 | Factual
no change in dimension of lump | 0 | 0 | Factual
multidisciplinary meeting | 0 | 0 | Factual
right mastectomy | 0 | 0 | Factual
axillary dissection | 0 | 0 | Factual
breast surgical wound healing regular | 24 | 24 | Factual
pathology assessment | 24 | 24 | Factual
fibroelastosis | 24 | 24 | Factual
chronic inflammation | 24 | 24 | Factual
isolated neoplastic cells | 24 | 24 | Factual
axillary nodes negative | 24 | 24 | Factual
restaging brain/chest/abdomen CT | 24 | 24 | Factual
no distant metastasis | 24 | 24 | Factual
BRCA and p53 mutation tests negative | 24 | 24 | Factual
autologous skin graft | 168 | 168 | Factual
no further complications | 168 | 168 | Factual
PICC implant | 168 | 168 | Factual
resumed chemotherapy | 168 | 0 | Factual
carboplatin | 168 | 0 | Factual
paclitaxel | 168 | 0 | Factual
dose reduction | 168 | 0 | Factual
good tolerance | 720 | 720 | Factual
completed fourth and last cycle | 720 | 720 | Factual
started follow-up | 720 | 720 | Factual