33 weeks gestation | 0
female | 0
vaginal delivery | 0
birth weight 1744 g | 0
Apgar score 9 at 1 minute | 0
Apgar score 9 at 5 minutes | 0
transfer to neonatal intensive care unit | 0
routine management of prematurity | 0
severe persistent hypoglycemia | 0
umbilical venous catheter placement | 48
maximum glucose infusion rate 21 mg/kg/min | 48
systolic murmur | 120
echocardiogram | 120
small patent ductus arteriosus | 120
umbilical venous catheter tip at foramen ovale | 120
removal of umbilical venous catheter | 120
fever | 168
tachypnea | 168
grunting | 168
thrombocytopenia | 168
platelets 81000 bil/L | 168
blood culture collection | 168
cerebrospinal fluid studies | 168
gentamicin initiation | 168
vancomycin initiation | 168
acyclovir initiation | 168
inadequate intravenous access | 168
persistent hypoglycemia | 168
need for antibiotics | 168
peripherally inserted central catheter attempted | 168
peripherally inserted central catheter failed | 168
bilious emesis episodes | 192
abdominal ultrasound negative | 192
upper gastrointestinal studies negative | 192
cranial ultrasound | 192
bilateral grade 1 intraventricular hemorrhages | 192
Broviac catheter insertion | 192
blood culture grew methicillin-sensitive Staphylococcus aureus | 192
cerebrospinal fluid no growth | 192
acyclovir discontinued | 192
cefotaxime added | 192
repeat echocardiogram | 240
5x5 mm mass in atrial septum | 240
Broviac pulled back | 240
mass persisted | 240
anticoagulation withheld | 240
repeat echocardiogram | 264
questionable increase in mass size | 264
gradual decrease in mass size | 264
no mass seen | 552
repeated cranial ultrasounds stable | 552
scalp nodule debrided | 408
leg nodule debrided | 408
methicillin-sensitive Staphylococcus aureus growth | 408
nafcillin course completed | 408
gentamicin course completed | 408
Broviac removed | 408
echocardiograms stable post-discharge | 408
no other sites of infection | 408
intra-atrial cardiac mass | 240
methicillin-sensitive Staphylococcus aureus | 192
conservative management | 240
