63 years old | 0
female | 0
admitted to the hospital | 0
general body malaise | -48
diarrhea | -48
vomiting | -48
influenza-like symptoms | -48
confusion | 0
splenectomy | -77496
idiopathic thrombocytopenic purpura | -77496
menometrorhagia | -77496
vaccinated with PPV23 | -672
fever | 0
hypotension | 0
bradycardia | 0
tachypnea | 0
decreased oxygen saturation | 0
cyanosis | 0
severe sepsis | 0
volume therapy | 0
broad-spectrum antimicrobial therapy | 0
hydrocortisone | 0
white blood cell count | 0
neutrophils | 0
hemoglobin | 0
thrombocytes | 0
C-reactive protein | 0
P-lactate | 0
aB-P-O2 | 0
aB-P-CO2 | 0
aB-pH | 0
Streptococcus pneumococcal urinary antigen test | 0
disseminated intravascular coagulation | 24
microthrombi | 24
blood cultures | 48
S. pneumoniae | 48
antimicrobial treatment | 48
penicillin G | 48
suspicion of endocarditis | 72
trans-thoracic echocardiography | 72
modest hypokinesia | 72
ejection fraction | 72
necrosis of the fingertips and toes | 72
renal insufficiency | 72
hemodialysis | 72
antibiotic therapy | 72
ceftriaxone | 72
leucocytes | 96
CRP | 96
fever | 96
tracheal secret | 96
culture | 96
transferred to the medical department | 216
antibiotics | 216
serological analysis | 216
pneumococcal isolate | 216
serotype 12F | 216
discharged | 528
oral dicloxacillin | 528
necrotic tissue | 528
wound cultures | 528
Staphylococcus aureus | 528
haemolytic streptococci group C/G | 528
amputated | 774
readmitted | 2160
severe sepsis | 2160
sepsis regimen | 2160
ceftriaxone | 2160
transesophageal echocardiography | 2160
endocarditis | 2160
aortic valve | 2160
blood cultures | 2160
S. pneumoniae | 2160
penicillin G | 2160
conservative treatment | 2160
recovered | 2448
antibody response | -77496
antibody response | -77496
antibody response | 0
antibody response | 528
antibody response | 2448