18 years old | 0
male | 0
admitted to the hospital | 0
backache | -30
calculi in both kidneys associated with ureteral calculi | -30
purulent urine | -30
severe fever | -30
chill | -30
low blood pressure | -30
blood and urine samples sent to the laboratory for culture | -30
empiric anti-infection drugs | -30
imipenem and Cilastatin sodium | -30
fluid resuscitation | -30
vasoactive agent (Norepinephrine) | -30
Hydrocortisone sodium succinate hormone | -30
anuric | -48
ARDS | -48
invasive ventilatory support with endotracheal intubation | -48
CRRT | -48
cold, clammy extremities | 0
loud bubbling sound in the lung | 0
arterial blood gas analysis | 0
oxygen partial pressure 50 mmHg | 0
lactic acid 10.6 mmol/L | 0
bicarbonate 10.8 mmol/L | 0
central venous pressure 20 cmH20 | 0
B lines in the lung | 0
cardiac function detected through the chest wall | 0
diffuse dysfunction, severe functional damage in the left ventricle | 0
LVEF 20.3% | 0
sinus tachycardia associated with broad ST depression | 0
elevated troponin I | 0
elevated amino-terminal brain natriuretic peptide precursor | 0
creatinine 356 μmol/L | 0
anuria | 0
ARDS | 0
sepsis-induced cardiomyopathy | 0
refractory septic shock | 0
VA-ECMO treatment initiated | 0
ECMO venous leading-out end used a 20F catheter | 0
ECMO arterial leading-in end used a 17F catheter | 0
arterial catheter placed in the right femoral artery | 0
ECMO ran normally 3000 rpm | 0
blood flow 3.5 L/min | 0
arterial pressure 135 mmHg | 0
venous pressure -29 mmHg | 0
Norepinephrine and Epinephrine stopped | 0.5
bedside CRRT performed | 0.5
lactic acid level declined | 2
vasoactive drugs stopped | 10
arterial blood lactate level reached the normal range | 12
extended-spectrum β-lactamase-positive Escherichia coli found in both blood and urine cultures | 48
inflammatory indices (e.g. leukocytes, calcitonin, C-reactive protein) decreased | 48
anti-infection regimen continued | 48
minimum serum trough concentration of Vancomycin monitored | 48
black and necrotic skin found at the extremities of both lower limbs and the end of a finger on the right upper limb | 120
patient successfully weaned from ECMO therapy | 144
renal function scaled as acute kidney injury grade 3 | 144
bedside CRRT discontinued | 144
patient began urinating | 144
vascular ultrasonography and computed tomography angiography performed in the bilateral lower limbs | 144
vascular surgery consultation | 144
necrotic tissues of the lower extremity amputated | 168
tracheal intubation | 168
spontaneous breathing successful | 168
trachea opened | 168
anti-infection combination of imipenem and Cilastatin sodium and Vancomycin replaced by Cefoperazone sodium and Sulbactam sodium | 168
bedside physical rehabilitation started | 168
patient weaned from the ventilator | 240
tracheotomy tube sealed | 252
patient discharged | 336
intermittent hemodialysis | 336
6-month follow-up | 336