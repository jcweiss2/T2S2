46 years old | 0
female | 0
admitted to the hospital | 0
multiple pelvic fractures | 0
multiple lacerations | 0
acute traumatic craniocerebral injury | 0
superficial skin contusion | 0
multiple burns | 0
debridement | 0
analgesics | 0
anti-infection | 0
hemostasis | 0
tetanus prevention | 0
wound exposure | 0
rehydration | 0
blood pressure dropped | 24
hemorrhagic shock | 24
intra-abdominal hemorrhage | 24
pelvic fracture | 24
transferred to ICU | 24
enhanced dilatation | 24
rehydration treatment | 24
anti-infection | 24
analgesia | 24
nutritional support | 24
single room isolation | 24
appropriate braking | 24
wound disinfection | 24
external application of burn cream | 24
exposure treatments | 24
intermittent moderate fever | 48
bilateral blood samples collected | 120
blood culture reports | 168
Pandoraea species isolated | 168
in vitro susceptibility testing | 168
antibiotic treatment changed | 216
imipenem | 216
tigecycline | 216
second blood culture reports | 240
Pandoraea species isolated | 240
bacteria culture | 288
high-throughput gene detection | 288
Pandoraea species isolated | 288
16S ribosomal RNA gene sequencing | 288
MALDI-TOF MS | 288
Pandoraea sputorum confirmed | 288
condition improved | 336
normal body temperature | 336
normal CRP | 336
normal PCT | 336
scanty wound exudation | 336
shifted to Department of Burn and Plastic Surgery | 336
wounds and fractures healed | 1440
discharged | 1440