67 years old | 0  
    woman | 0  
    right-sided headaches | -2928  
    visual disturbance | -2928  
    acute confusion | -720  
    fever | -720  
    vomiting | -720  
    photophobia | -720  
    right-sided radicular leg pain | -720  
    extreme lethargy | -720  
    thirst | -720  
    weight loss | -720  
    loss of appetite | -720  
    new onset nocturia | -720  
    hyponatraemia | -720  
    primary breast carcinoma | -8760  
    Grade 2 tumor | -8760  
    ER+ | -8760  
    PR+ | -8760  
    HER2* | -8760  
    lymph node negative | -8760  
    wide local excision | -8760  
    post-operative radiotherapy | -8760  
    letrozole | -8760  
    brain MRI | -2880  
    partly solid tumor | -2880  
    partly cystic suprasellar tumor | -2880  
    compression of optic apparatus | -2880  
    repeat MRI | -2880  
    progression of tumor | -2880  
    widespread metastatic lesions | -2880  
    MRI spine | -720  
    intradural extramedullary lesion | -720  
    equivocal pial nodules | -720  
    radiological diagnosis of craniopharyngioma | 0  
    rapid increase in size | 0  
    differential diagnosis of breast metastasis | 0  
    differential diagnosis of hypothalamic glioma | 0  
    no visceral metastatic disease | 0  
    CT chest | 0  
    CT abdomen | 0  
    CT pelvis | 0  
    multidisciplinary team meeting | 0  
    stealth-guided endoscopic resection | 0  
    CSF cytology | 0  
    lumbar puncture | 0  
    intraoperative smear | 0  
    histology | 0  
    squamous epithelial cells | 0  
    moderate pleomorphism | 0  
    focal keratinisation | 0  
    granulation tissue | 0  
    chronic lymphocytic inflammation | 0  
    cytokeratins positive (MNF116, CK7, CK5/6) | 0  
    CK20 negative | 0  
    TTF1 negative | 0  
    scattered cells within granulation tissue | 0  
    increased Ki-67 proliferation | 0  
    molecular sequencing BRAF V600K mutation | 0  
    lumbar puncture 4 weeks post-surgery | 672  
    squamous cells compatible with papillary craniopharyngioma | 672  
    pancytokeratin positive | 672  
    CK7 positive | 672  
    EMA positive | 672  
    GATA3 negative | 672  
    GCDFP-15 negative | 672  
    ER negative | 672  
    PR negative | 672  
    BRAF V600K mutation in CSF | 672  
    atypical squamous epithelial cells in CSF | 672  
    CSF seeding | 672  
    metastatic deposits | 672  
    malignancy confirmed | 672  
    Ki67 index elevated | 672  
    inflammatory response | 672  
    BRAF inhibitors considered | 672  

