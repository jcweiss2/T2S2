24 years old | 0
female | 0
pregnant | 0
admitted to the hospital | 0
abdominal pain | -120
abdominal distension | -120
constipation | -120
diagnosed with preterm delivery | -120
evaluated by surgical and obstetric teams | 0
dehydrated | 0
hypotension | 0
tachycardia | 0
tachypnea | 0
asymmetrically distended abdomen | 0
tenderness all over abdomen | 0
rectum empty on digital examination | 0
foetal viability assessed | 0
vaginal examination not suggestive of threatened preterm labour | 0
elevated white cell count | 0
urine analysis clear | 0
ultrasound scan of abdomen and pelvis | 0
distended bowel loop | 0
moderate amount of free fluid in peritoneal cavity | 0
single viable foetus | 0
clinical diagnosis of IO proposed | 0
abdominal X-ray | 0
dilated large bowel | 0
abnormal gas pattern | 0
coffee bean appearance | 0
sigmoid volvulus diagnosed | 0
gastroenterology team consulted | 0
emergency sigmoidoscopy | 0
twisted sigmoid colon confirmed | 0
obstruction not negotiable | 0
foetal distress | 0
deceleration in heart rate | 0
concomitant caesarean section decided | 0
premature foetus delivered | 24
male preterm infant | 24
weight 750g | 24
admitted to neonatal ICU | 24
mechanical ventilation | 24
gangrenous sigmoid colon | 24
necrosis | 24
sigmoid mesocolon twisted | 24
necrotic colon posteriorly displaced | 24
lower segment caesarean section | 24
Hartmann’s procedure | 24
end colostomy fashioned | 24
rectal stump closed | 24
post-operative course uneventful | 24
discharged home | 216
child discharged home | 720
reversal of Hartmann’s | 2160
bowel continuity restored | 2160
colo-rectal anastomosis | 2160