2 years old | 0
male | 0
domestic shorthair cat | 0
castrated | 0
admitted to the hospital | 0
progressive signs of weakness | 0
neurologic dysfunction | 0
history of chronic kidney disease | -672
leukocytosis | -2
neutrophilia | -2
lymphocytosis | -2
mild azotemia | -2
blood urea nitrogen | -2
creatinine | -2
ataxia | -2
vomiting | -2
tetraparesis | -2
bradycardia | 0
tachypnea | 0
stuporous mentation | 0
tetraplegia | 0
absent withdrawals | 0
absent peripheral reflexes | 0
weak gag reflex | 0
absent menace | 0
short shallow breaths | 0
mild hypercapnia | 0
mild azotemia | 0
baclofen ingestion | -4
ingestion of 10 mg baclofen tablet | -4
hemodialysis | 1.5
IV fluid therapy | 1.5
lactated Ringer’s solution | 1.5
hemodialysis catheter placement | 1.5
mechanical ventilation | 2
propofol administration | 2
endotracheal intubation | 2
manual ventilation | 2
severe hemorrhage | 2
hypotension | 2
tachycardia | 2
heparin therapy discontinuation | 2
hypertonic saline administration | 2
packed RBCs administration | 2
fresh frozen plasma administration | 2
heparin therapy restart | 2
hemodialysis completion | 5
weaning from ventilator | 5
extubation | 5
improvement in muscle tone | 6
weakly ambulatory | 6
resolution of hypercapnia | 7
resolution of acidemia | 7
complete resolution of neurologic signs | 12
discharge | 24
follow-up appointment | 168
normal behavior | 168
normal appetite | 168
persistent mild azotemia | 168
non-regenerative anemia | 168
aggregate reticulocyte count | 168
normal white blood cell count | 168
continuing treatment for CKD | 720
doing well | 720