57 years old | 0  
    male | 0  
    admitted for unrelated peripheral blood stem cell transplantation | 0  
    Philadelphia-positive acute lymphoblastic leukemia | -1440  
    remission-induction chemotherapy | -1440  
    five cycles of intrathecal chemotherapy | -1440  
    pre-transplant conditioning chemotherapy with fludarabine | -216  
    melphalan | -216  
    anti-thymocyte immunoglobulin | -216  
    ciprofloxacin prophylaxis | -216  
    itraconazole syrup prophylaxis | -216  
    acyclovir prophylaxis | -216  
    stem cell transplantation | -48  
    neutropenia developed | -48  
    neutropenia progressed | -48  
    intermittent mild abdominal pain | -96  
    diarrhea | -96  
    chronic diarrhea before hospitalization | -216  
    Clostridium difficile toxin assay | -216  
    culture done at hospital day 5 | -216  
    severe pain at left chest wall, left buttock, and thigh | 0  
    localized swelling | 0  
    tissue edema progressed rapidly | 0  
    no obvious traumatic injury | 0  
    intravenous Hickman catheter | 0  
    no infectious signs at exit site | 0  
    empirical antibiotics started with piperacillin/tazobactam | 0  
    vancomycin started | 0  
    hemoglobin 9.3 g/dL | 0  
    hematocrit 25.2% | 0  
    white blood cells 10/mm3 | 0  
    absolute neutrophil count 0/mm3 | 0  
    platelet 61,000/mm3 | 0  
    ciprofloxacin discontinued | 0  
    chest X-ray showed soft tissue swelling with air density | 0  
    blood pressure fell to 92/60 mmHg | 0  
    heart rate 164/min | 0  
    oxygen saturation 83% | 0  
    normal saline administration | 0  
    oxygen applied via simple facial mask | 0  
    vital signs stabilized | 0  
    chest and abdominal computed tomography revealed multiple emphysematous soft tissue infections | 0  
    needle aspiration from soft tissue lesion | 0  
    heart rate increased to 163/min | 10  
    blood pressure 98/63 mmHg | 10  
    planned transfer to intensive care unit | 10  
    cardiac arrest occurred | 12  
    cardiopulmonary resuscitation | 12  
    death without return of spontaneous circulation | 12  
    Clostridium perfringens isolated from blood cultures | 12  
    Clostridium perfringens isolated from aspirated fluid culture | 12  

    57 years old | 0
male | 0
admitted for unrelated peripheral blood stem cell transplantation | 0
Philadelphia-positive acute lymphoblastic leukemia | -1440
remissionEinduced chemotherapy | -1440
five cycles of intrathecal chemotherapy | -1440
preEtransplant conditioning chemotherapy with fludarabine | -216
melphalan | -216
antiEthymocyte immunoglobulin | -216
ciprofloxacin prophylaxis | -216
itraconazole syrup prophylaxis | -216
acyclovir prophylaxis | -216
stem cell transplantation | -48
neutropenia developed | -48
neutropenia progressed | -48
intermittent mild abdominal pain | -96
diarrhea | -96
chronic diarrhea before hospitalization | -216
Clostridium difficile toxin assay | -216
culture done at hospital day 5 | -216
severe pain at left chest wall, left buttock, and thigh | 0
localized swelling | 0
tissue edema progressed rapidly | 0
no obvious traumatic injury | 0
intravenous Hickman catheter | 0
no infectious signs at exit site | 0
empirical antibiotics started with piperacillin/tazobactam | 0
vancomycin started | 0
hemoglobin 9.3 g/dL | 0
hematocrit 25.2% | 0
white blood cells 10/mm3 | 0
absolute neutrophil count 0/mm3 | 0
platelet 61,000/mm3 | 0
ciprofloxacin discontinued | 0
chest XEray showed soft tissue swelling with air density | 0
blood pressure fell to 92/60 mmHg | 0
heart rate 164/min | 0
oxygen saturation 83% | 0
normal saline administration |0
oxygen applied via simple facial mask |0
vital signs stabilized |0
chest and abdominal computed tomography revealed multiple emphysematous soft tissue infections |0
needle aspiration from soft tissue lesion |0
heart rate increased to 163/min |10
blood pressure 98/63 mmHg |10
planned transfer to intensive care unit |10
cardiac arrest occurred |12
cardiopulmonary resuscitation |12
death without return of spontaneous circulation |12
Clostridium perfringens isolated from blood cultures |12
Clostridium perfringens isolated from aspirated fluid culture |12