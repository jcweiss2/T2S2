29 years old | 0
male | 0
African American | 0
admitted to the hospital | 0
sickle cell disease | -8760
hemosiderosis | -8760
cirrhosis | -8760
vaso-occlusive pain crisis | 0
uncontrolled epistaxis | 0
deferasirox | -8760
folic acid | -8760
oxycodone | -8760
denies tobacco | 0
denies alcohol | 0
denies drug use | 0
jaundiced | 0
alert | 0
fully oriented | 0
abdomen soft | 0
no tenderness | 0
no organomegaly | 0
normal bowel sounds | 0
new-onset confusion | 24
hepatic encephalopathy | 24
conjugated hyperbilirubinemia | 0
total serum bilirubin 57 mg/dL | 0
direct serum bilirubin 30 mg/dL | 0
alkaline phosphatase 306 U/L | 0
aspartate transaminase 227 U/L | 0
alanine transaminase 54 U/L | 0
white blood cell count 38.6 k/µL | 0
hemoglobin 6.3 g/dL | 0
platelet count 39 k/µL | 0
Coomb's testing negative | 0
fibrinogen 412 mg/dL | 0
INR 2.3 | 0
model for end-stage liver disease-sodium score 40 | 0
acute kidney injury | 0
serum creatinine 3.48 mg/dL | 0
cirrhotic liver morphology | 0
patent hepatic vasculature | 0
appropriate flow | 0
changes consistent with cirrhosis | 0
no biliary ductal dilatation | 0
acute-on-chronic liver failure | 0
multi-system organ failure | 0
acute sickle cell intrahepatic cholestasis | 0
intubation | 0
mechanical ventilation | 0
acute hypoxic respiratory failure | 0
acute chest syndrome | 0
vancomycin | 0
meropenem | 0
exchange transfusion | 0
HbS level 56.3 g/dL | 0
HbS level 8.2 g/dL | 0
hepatic synthetic function did not improve | 0
listed for liver transplantation | 0
model for end-stage liver disease-sodium score 40 | 0
liver transplantation | 216
HCV NAT positive donor | 216
HCV NAT negative patient | 216
glecaprevir/pibrentasvir | 239
sustained virologic response | 744
tacrolimus | 216
mycophenolate mofetil | 216
steroid taper | 216
immunosuppression induction therapy | 216
antithymocyte globulin | 216
HCV ribonucleic acid > 100000000 IU/mL | 72
HCV genotype 1A | 72
exchange transfusion resumed | 216
monthly exchange transfusions | 744
target HbS < 20% | 744
liver synthetic function preserved | 8760
chronic tacrolimus immune suppressive therapy | 8760