40 years old | 0
male | 0
admitted to the hospital | 0
fever | -96
nausea | -96
vomiting | -96
enlarging non-tender left neck swelling | -96
hypotensive | 0
febrile | 0
confused | 0
unilateral anterior cervical triangle swelling | 0
erythematous rash | 0
left side of neck | 0
anterior chest wall | 0
sinus rhythm | 0
left anterior fascicular block | 0
intravenous fluid resuscitation | 0
broad-spectrum antibiotics | 0
elevated inflammatory markers | 0
C-reactive protein 205 mg/L | 0
computed tomography neck and thorax | 0
acute inflammatory process | 0
left submandibular space | 0
unilateral enlarged lymph nodes | 0
necrotizing lymphadenopathy | 0
septic shock | 24
normal haemoglobin | 24
neutrophils | 24
elevated inflammatory markers | 24
lymphopoenia | 24
thrombocytopoenia | 24
hyponatraemia | 24
hepatitis | 24
hypoalbuminaemia | 24
coagulopathy | 24
myocarditis | 24
troponin T 1104 ng/L | 24
NT-proBNP 48 412 pg/mL | 24
viral and bacterial investigations | 24
negative | 24
vasculitis screen | 24
negative | 24
transthoracic echocardiogram | 24
normal left ventricular function | 24
moderate central mitral regurgitation | 24
ultrasound-guided biopsy | 72
left anterior cervical lymph node | 72
suppurative necrotizing lymphadenitis | 72
new erythema of the oral mucosa | 96
fissured lips | 96
strawberry tongue | 96
bilateral conjunctival injection | 96
intravenous immunoglobulins | 96
high-dose aspirin | 96
dramatic clinical improvement | 120
acute transient left upper limb weakness | 240
CT angiogram | 240
magnetic resonance imaging | 240
vertebral artery dissection | 240
negative | 240
stroke | 240
negative | 240
computed tomography coronary angiography | 720
cardiac magnetic resonance imaging | 720
two sequential aneurysms | 720
right coronary artery | 720
left anterior descending artery | 720
no associated thrombus | 720
mural thickening | 720
coronary plaque | 720
perivascular fatty changes | 720
normal left ventricular volumes | 720
preserved function | 720
focal regions of mid-wall fibrosis | 720
previous myocarditis | 720
follow-up CTCA | 2880
resolution of the LAD aneurysm | 2880
improvement of the two focal aneurysms | 2880
right coronary artery | 2880
discharged | 240