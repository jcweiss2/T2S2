36 years old | 0
Hispanic | 0
gravida 3 | 0
para 0 | 0
17 weeks' gestation | 0
lower abdominal pain | -48
mild complaints | -24
discharged home | -24
diagnosis of intestinal gas | -24
persistent pain | 0
severe pain | 0
exacerbated by movement | 0
loss of appetite | 0
no nausea | 0
no emesis | 0
tachycardic | 0
involuntary guarding | 0
suprapubic region | 0
sterile speculum examination | 0
normal closed cervix | 0
spontaneous rupture of yellow purulent fluid | 0
posterior vaginal fornix | 0
posterior vaginal wall defect | 0
elevated white blood cell count | 0
neutrophilic shift | 0
transvaginal ultrasound | 0
complex collection in posterior cul-de-sac | 0
multiloculated abscess | 0
pelvic magnetic resonance imaging | 0
right ovarian torsion | 0
abscess formation | 0
antibiotic treatment | 0
ceftriaxone | 0
metronidazole | 0
general surgery team consulted | 0
sepsis | 24
worsening hypotension | 24
pain | 24
multidisciplinary meeting | 24
vancomycin | 24
operating room | 24
diagnostic laparoscopy | 24
general surgery team | 24
obstetrics/gynecology team | 24
examination under anesthesia | 24
defect in posterior fornix | 24
purulent fluid | 24
appendix adherent to uterus | 24
abscess | 24
right fallopian tube | 24
right ovary | 24
adhesions | 24
right lower quadrant | 24
Penrose drain | 24
fetal status | 24
reassuring | 24
postoperative day 5 | 120
piperacillin–tazobactam | 120
regular diet | 120
Penrose drain removal | 120
discharged | 120
oral cefpodoxime | 120
recovery | 120
office follow-up visit | 168
uncomplicated normal spontaneous vaginal delivery | 2808
401/7 weeks | 2808
healthy infant | 2808
no malformations | 2808
no neurological sequelae | 2808
no behavioral sequelae | 2808
appendicitis | -48
peritoneovaginal fistula | 24
isolated appendiceal endometriosis | 24
decidualization | 24
endometriosis | 24
acute inflammatory infiltrates | 24
neutrophils | 24
appendiceal endometriosis | 24
perforation | 24
peritonitis | 24
abscess development | 24
inflammatory response | 24
decidua | 24
endometriotic appendix | 24