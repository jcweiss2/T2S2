39 years old | 0
female | 0
admitted to the hospital | 0
sepsis | 0
piperacillin-tazobactam | 0
renal cell carcinoma | -1560
left partial nephrectomy | -1560
interferon | -936
bevacizumab | -936
shortness of breath | 12
tachypnea | 12
chest discomfort | 12
decreased breath sounds | 12
tympanic percussion | 12
trachea deviation | 12
bilateral jugular stasis | 12
low saturation | 12
oxygen therapy | 12
thoracocentesis | 12
air escape | 12
hydropneumothorax | 12
contralateral mediastinal shift | 12
chest drain | 12
turbid brownish fluid | 12
non-invasive mechanical ventilation | 24
chest discomfort improved | 48
lung expansion | 48
nasogastric feed | 48
pleural effusion | 48
neutrophilic exudate | 48
low pH | 48
low protein | 48
normal glucose | 48
high lactate dehydrogenase | 48
high amylase | 48
esophageal perforation suspected | 48
methylene blue test | 72
gastropleural fistula | 72
computed tomography | 72
parenteral nutrition | 96
sudden bleeding | 120
hypovolemic shock | 120
fluid resuscitation | 120
blood transfusion | 120
vasopressor support | 120
upper gastrointestinal endoscopy | 120
blood clot | 120
embolization of splenic arteries | 144
no further bleeding | 144
palliative care | 168
death | 240
shock | 240
acute respiratory insufficiency | 240