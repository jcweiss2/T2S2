30 years old | 0
male | 0
idiopathic bronchiectasis | 0
admitted to the emergency department | 0
fever | 0
productive cough | 0
chest pain | 0
dyspnea | 0
anosmia | 0
contact with recovered COVID-19 friend | -72
bilateral crackles at lower lobes | 0
peripheral oxygen saturation 65% | 0
no respiratory distress | 0
connected to high flow nasal cannula | 0
chest X-ray showing peripheral infiltrates | 0
desaturated SpO2 55% | 0
intubated | 0
mechanical ventilation | 0
COVID-19 confirmed by RT-PCR | 0
normal electrocardiogram | 0
normal cardiac enzymes | 0
normal echocardiography | 0
leukocytosis 17.9×10⁹/L | 0
lymphocytopenia 0.42×10⁹/L | 0
increased D-dimer 3.3 mcg/ml | 0
increased C-reactive protein 245 mg/liter | 0
increased lactate dehydrogenase 904 units/liter | 0
increased ferritin 883 ng/ml | 0
contrast chest CT scans excluded pulmonary embolism | 0
bilateral peripheral ground-glass opacities | 0
bronchiectasis on CT | 0
admitted to COVIDE-19 ICU | 0
diagnostic work-up for infections | 0
serum 25(OH)D levels measured | 0
lockdown for three months | -2160
empiric therapy with ribavirin | 0
empiric therapy with ceftriaxone | 0
empiric therapy with azithromycin | 0
prophylactic anticoagulation | 0
ARDS-net ventilation | 0
prone position ventilation | 0
supportive ICU care | 0
no improvement in respiratory status on day-3 | 72
Bordetella bronchiseptica culture ≥105 cfu/ml | -24
antibiotic regime adjusted | 72
doxycycline received for two weeks | 72
severe vitamin D deficiency 25 nmol/L | 0
vitamin D3 bolus 100,000 IU | 72
weekly vitamin D3 25,000 IU | 72
extubated on day-15 | 360
RT-PCR negative for COVID-19 on day-18 | 432
microbiology negative on day-18 | 432
discharged on day-20 | 480
monitor pet dog for kennel cough | 480
review vitamin D supplementation | 480
review dietary habits | 480
happy hypoxemia | 0
cytokine storm | 0
Bordetella bronchiseptica infection | -24
fulminant clinical presentation | 0
vitamin D deficiency linked to severity | 0
combination therapy improvement | 0
no known competing interests | 0
admitted to COVID-19 ICU | 0
prone position ventilation |&nbsp;0
