throat pain | -168
odynophagia | -168
blood tests | -168
diagnosis of acute promyelocytic leukemia | -168
treatment with daunorubicin plus vesanoid | -168
physical examination | 0
necrotic lesion in the M. palatoglossus, soft palate, uvula and right tonsil | 0
unpleasant odor | 0
biopsy | 0
culture | 0
histopathologic findings showed nonspecific chronic diffuse inflammation | 0
necrotic areas and numerous bacteria | 0
culture identified Enterococcus spp, Staphylococcus aureus and Candida SP | 0
diagnosis of noma-like lesion | 0
antibiotic therapy using ceftazidime, amicacin, vancomycin, fluconazole and penicillin G | 0
pneumonia | 24
sepsis | 24
treatment in the intensive care unit | 24
total recovery | 45
extensive loss of soft palate tissue | 45
measles | -10000
rubella | -10000
typhoid fever | -10000
whooping cough | -10000
typhus | -10000
syphilis | -10000
tuberculosis | -10000
leukemia | -10000
mucocutaneous leishmaniasis | -10000
lupus erythematosus | -10000
leprosy | -10000
agranulocytic ulcerations | -10000
physical trauma | -10000
oral cancer | -10000
yaws | -10000 
no shortness of breath | 0
denies chest pain | 0