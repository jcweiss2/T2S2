57 years old | 0
male | 0
dyspnea | -48
cough | -48
sputum | -48
left shoulder pain | -48
diaphoresis | -48
myalgia | -48
fever | -48
chilled sensation | -48
diabetes mellitus | -2628
smoker | -2628
alcohol consumption | -2628
exposure to marble dust | -2628
linagliptin | -2628
metformin | -2628
admitted to the hospital | 0
blood pressure 206/109 | 0
heart rate 123 beats/minute | 0
body temperature 38.2°C | 0
left hydropneumothorax | 0
pleural adhesion | 0
leukocytosis | 0
erythrocyte sedimentation rate 121 mm/hr | 0
C-reactive protein level 45.8 mg/dL | 0
arterial partial pressure of oxygen 50.9 mmHg | 0
oxygen therapy | 0
hemoglobin A1c level 6.9% | 0
aspartate aminotransferase 21 IU/L | 0
alanine aminotransferase 26 IU/L | 0
total bilirubin 0.5 mg/dL | 0
prothrombin time 1.18 INR | 0
albumin concentration 3.0 g/dL | 0
blood cultures | 0
pleural fluid sample | 0
turbid pleural fluid | 0
thick pleural fluid | 0
brownish-yellow pleural fluid | 0
foul odor | 0
exudative pleural fluid | 0
intravenous ceftriaxone | 0
intravenous levofloxacin | 0
intravenous clindamycin | 0
24-French chest tube insertion | 0
admitted to intensive care unit | 0
esophago-gastro-duodenoscopy | 24
no esophageal injury | 24
micro-rupture possibility | 24
culture results | 120
K. kristinae identification | 120
antibiotic treatment escalation | 216
intravenous piperacillin-tazobactam | 216
intravenous levofloxacin | 216
relapsed fever | 216
discharged | 552
amoxicillin-clavulanic acid prescription | 552
follow-up blood culture negative | 240
improved chest radiographic findings | 552