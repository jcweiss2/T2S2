54 years old | 0
    male | 0
    presented following motor vehicle collision | 0
    Glasgow Coma Scale 13 | 0
    Glasgow Coma Scale declined | 0
    intubated | 0
    admitted to surgical ICU | 0
    C1 transverse foramen fracture | 0
    bilateral rib fractures | 0
    pulmonary contusions | 0
    became febrile shortly after admission | 24
    lower respiratory culture consistent with polymicrobial pneumonia | 0
    started on broad-spectrum antibiotics | 0
    family provided history of active crack cocaine use | 48
    restarted on quetiapine 400 mg at bedtime | 48
    restarted on mirtazapine 30 mg at bedtime | 48
    persistent intermittent agitation | 48
    agitation difficult to control despite opioids | 48
    agitation difficult to control despite dexmedetomidine | 48
    agitation difficult to control despite lorazepam | 48
    received intravenous haloperidol 5 mg for agitation | 120
    febrile to 102.2°F–104.7°F | 144
    acetaminophen | 144
    cooling blanket | 144
    ice saline gastric lavage | 144
    developed tachycardia | 144
    developed hypertension | 144
    diffuse lead-pipe rigidity | 144
    hyperreflexia | 144
    two-beat clonus | 144
    differential diagnosis broadened to include sepsis | 144
    differential diagnosis broadened to include NMS | 144
    differential diagnosis broadened to include serotonin syndrome | 144
    differential diagnosis broadened to include cocaine withdrawal | 144
    serum creatine kinase 247 IU/L | 144
    received IV dantrolene 2.5 mg/kg | 144
    quetiapine discontinued | 144
    mirtazapine discontinued | 144
    haloperidol discontinued | 144
    dysautonomia resolved | 144.5
    rigidity resolved | 144.5
    hyperreflexia resolved | 144.5
    temperature downtrended | 144.5
    blood cultures sent | 144
    urine cultures sent | 144
    lower respiratory cultures sent | 144
    continued on maintenance oral dantrolene | 168
    resolution of rigidity | 168
    improvement in fever curve | 168
    bromocriptine added | 192
    dantrolene discontinued | 240
    rigidity recurred | 264
    hyperreflexia recurred | 264
    dantrolene restarted | 264
    tapered 14-day course | 264
    passed spontaneous breathing trial | 312
    extubated | 312
    mental status returned to baseline | 312
    no further recurrence of symptoms | 312
    resumed quetiapine 50 mg QHS | 528
    discharged | 696
    no shortness of breath | 0
    denies chest pain | 0
    