46 years old | 0
man | 0
obesity | 0
body mass index 42 kg/m2 | 0
presented to emergency department | 0
right lower extremity weakness | -24
nausea | -24
generalized weakness | -24
diagnosed with SARS-CoV-2 infection | -1440
mild flu-like symptoms | -1440
positive total antibodies | -1440
two negative nasopharyngeal polymerase chain reaction | -1440
admission | 0
alert | 0
oriented | 0
hypotensive | 0
blood pressure 88/37 mmHg | 0
hypoxic | 0
oxygen saturation 89% | 0
nasal cannula at 3 L/min | 0
bilateral rhonchi | 0
right lower extremity strength 3/5 | 0
no skin rashes | 0
negative nasopharyngeal PCR | 0
positive total antibody test | 0
SARS-CoV-2 total antibodies 238 s/co ratio | 0
IgG 11 s/co ratio | 0
ferritin 962 ng/mL | 0
IL-6 121.09 pg/mL | 0
CRP 2.9 mg/dL | 0
LDH 802 units/L | 0
procalcitonin 0.678 ng/mL | 0
acute kidney injury | 0
creatinine 4.10 mg/dL | 0
high anion gap metabolic acidosis | 0
lactic acidosis | 0
chest x-ray left retrocardiac opacity | 0
no evidence of overt edema | 0
EKG NSTEMI | 0
troponin 0.282 ng/mL | 0
BNP 3590 pg/mL | 0
transthoracic echocardiography normal ejection fraction | 0
borderline elevated RVSP | 0
CT chest dependent ground glass opacities | 0
CT abdomen hepatic steatosis | 0
concern for posterior circulation stroke | 0
right ataxia | 0
mild right hemiparesis | 0
left hemianesthesia | 0
CT head unremarkable | 0
hypoxia | 0
required oxygen support 6 L nasal cannula | 0
hospitalization day 1 | 24
chest x-ray diffuse bilateral opacities | 24
tachypneic | 24
worsening hypoxemia | 24
required 40 L/min high-flow nasal cannula | 24
transferred to ICU | 24
invasive mechanical ventilation | 24
norepinephrine | 24
ceftriaxone 2 gm daily | 24
azithromycin 500 mg daily | 24
dexamethasone 6 mg daily | 24
unfractionated heparin | 24
repeat nasopharyngeal PCR negative | 24
hospitalization day 3 | 72
BAL PCR negative | 72
consultation with CDC | 72
high suspicion for MIS-A | 72
treated with tocilizumab 8 mg/kg | 72
steroids | 72
troponin 2.1 ng/mL | 72
BNP 5940 pg/mL | 72
repeat TTE RVSP 39.4 mmHg | 72
normal left ventricle | 72
normal left ventricular wall thickness | 72
normal left ventricular wall motion | 72
normal right ventricle | 72
kidney function deterioration | 72
CVVH | 72
hospitalization day 4 | 96
hospitalization day 5 | 120
no clinical improvement | 120
ferritin 1993 ng/mL | 120
IL-6 1412.44 pg/mL | 120
LDH 4773 units/L | 120
d-dimer 0.62 mcg/mL | 120
CRP 8.3 mg/dL | 120
liver function worsening | 120
kidney function worsening | 120
troponin persistently elevated | 120
multiorgan failure | 120
hospitalization day 6 | 144
requiring less ventilator support | 144
no pressors needed | 144
hospitalization day 8 | 192
hypotensive | 192
febrile | 192
thick foul-smelling respiratory secretions | 192
respiratory cultures Candida albicans | 192
vancomycin | 192
cefepime | 192
norepinephrine restarted | 192
ferritin >100,000 ng/mL | 192
LDH >12,000 units/L | 192
repeat SARS-CoV-2 PCR negative | 192
whole genome sequencing failed | 192
hospitalization day 9 | 216
hydrocortisone 50 mg q6h | 216
severe refractory acidosis | 216
hyperkalemia | 216
arrhythmia | 240
death | 240
negative respiratory viral panel | 0
negative HIV | 0
negative hepatitis C | 0
negative influenza | 0
no splenomegaly | 0
no cytopenia | 0
no hypofibrinogenemia | 0
no pericarditis | 0
no acute infarctions | 0
no skin lesions | 0
no malignancy | 0
no pulmonary embolism | 0
no vasculitis | 0
no sHLH | 0
no cytokine storm | 0
no re-infection | 0
negative BAL PCR | 72
negative BAL sequencing | 192
no IVIG administered | 0
no anakinra administered | 0
no additional tocilizumab doses | 0
no clinical trials | 0
funding none | 0
no conflict of interest | 0
