22 years old | 0
female | 0
admitted with abdominal distention | 0
vomiting | -168
constipation | -168
hyperventilation episodes | -168
Rett syndrome diagnosis | -173328
seizure disorders | -173328
air swallowing | -173328
difficulty in evacuation of stool | -173328
use of rectal enema | -173328
rectal digitation for defecation | -173328
no stool discharge for 4 days | -168
abdominal distension | 0
abdominal tenderness | 0
rebound | 0
septic appearance | 0
bloody discharge in rectal examination | 0
increased sphincter tonus | 0
decreased Turgol-tonus | 0
dilated bowel segments on X-ray | 0
air-fluid levels on X-ray | 0
coffee-bean sign on lower left quadrant | 0
acute abdomen due to sigmoid volvulus | 0
normal coagulation function | 0
normal liver function | 0
increased Blood Urea Nitrogen | 0
increased creatinine | 0
increased white blood cell count | 0
increased serum sodium | 0
increased blood glucose | 0
increased plasma CRP levels | 0
acute metabolic acidosis | 0
sinus tachycardia | 0
QT interval 500 ms | 0
urgent laparotomy | 0
sigmoid volvulus | 0
2 cm hard mass resembling colon tumor | 0
several hard nodular lesions in the liver | 0
Hartman procedure | 0
liver biopsy | 0
followed with septic shock | 24
intensive care management | 24
deteriorated pulmonary function | 24
deteriorated cardiac function | 24
death | 48
musinous adenocarcinoma (3 cm) | 48
liver metastasis adenocarcinoma | 48
no genetic analysis performed | 48
chronic constipation | -173328
swallowing problems | -173328
emergency operation due to gastrointestinal pathologies | 0
late hospital admission | -168
decreased pain sensation | -173328
septic shock complication | 24
colon cancer | 0
liver metastasis | 0
MECP2 gene mutation | -173328
hypermethylation of tumor suppressor genes | 48
scoliosis | 0
