12 years old | 0
female | 0
admitted to the burn center | 0
deep burns | 0
burns in 46% of total body surface area | 0
serial excision and grafting | 0
treated with broad-spectrum antibiotics | 0
severe sepsis | 0
complained of pain | 552
decreased visual acuity | 552
ophthalmologic examination | 552
best corrected visual acuity (BCVA) was hand motion in the right eye | 552
best corrected visual acuity (BCVA) was 20/20 in the left eye | 552
panuveitis | 552
anterior chamber hypopyon | 552
dense vitritis | 552
large chorioretinal abscess | 552
smear and culture of the vitreous biopsy | 552
Candida albicans | 552
diagnosed with fungal endogenous endophthalmitis | 552
treated with systemic fluconazole | 552
intravitreal injection of Amphotericin B | 552
pars plana deep vitrectomy | 552
BCVA was hand motion in the right eye | 1240
large macular scar | 1240
free from inflammation | 1240
left eye was normal | 1240
retinal detachment | 1488
repeat pars plana vitrectomy | 1488
membrane peeling | 1488
silicone oil injection | 1488
final BCVA improved to counting fingers (CF) at two meters | 2208
retina was completely attached | 2208
central macular scar | 2208