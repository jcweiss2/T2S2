22 years old | 0
female | 0
distant history of alcohol use | -672
distant history of cocaine use | -672
nausea | -168
vomiting | -168
subjective fevers | -168
myalgias | -168
fatigue | -168
denies chest pain | 0
denies dyspnea | 0
denies cough | 0
sinus tachycardia | 0
temperature of 36.9 degrees Celsius | 0
blood pressure of 75/40 mmHg | 0
oxygen saturations of 90% on room air | 0
elevated jugular venous pressure | 0
heart sounds difficult to hear on auscultation | 0
elevated white blood cell count | 0
neutrophil count of 13.0 × 10^9/L | 0
normal cardiac troponin I | 0
normal creatinine | 0
normal electrolytes | 0
normal beta-HCG | 0
negative urine toxicology | 0
sinus tachycardia with small voltages in the limb leads on ECG | 0
generous sized cardiac silhouette on chest X-ray | 0
clear lung fields on chest X-ray | 0
admitted to intensive care unit | 0
given fluids | 0
given ionotropic support with norepherine | 0
pipericillin-tazobactam started | 0
vancomycin started | 0
nasopharyngeal swab conducted | 0
nasopharyngeal swab positive for Influenza A H1N1 | 0
oseltamivir initiated | 0
remained hypotensive | 0
echocardiogram performed | 12
moderate sized pericardial effusion | 12
maximal diameter of 1.5 cm in maximal width | 12
right ventricular diastolic collapse | 12
significant respiratory variation seen on mitral valve annular doppler velocity | 12
urgent pericardiocentesis conducted | 12
immediate improvement of hemodynamic status | 12
withdrawal of all ionotropic support | 12
pericardial drain inserted | 12
repeat echocardiogram conducted | 48
resolution of pericardial effusion | 48
absence of echocardiographic findings of tamponade | 48
pericardial effusion negative for bacterial cultures | 48
pericardial effusion negative for acid fast bacilli | 48
pericardial effusion negative for malignancy | 48
serologic testing for HIV negative | 48
serologic testing for Hepatitis B negative | 48
serologic testing for Hepatitis C negative | 48
high dose ibuprofen initiated | 48
colchcine initiated | 48
pericardial drain removed | 120
repeat echocardiogram conducted | 168
no return of pericardial effusion | 168
discharged from hospital | 168