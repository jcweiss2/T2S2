61 years old | 0
male | 0
diabetic | 0
admitted to the emergency department | 0
generalized worsening | -168
fever | -168
dysphagia | -168
cervical swelling | -168
impacted fish bones in throat | -168
examined by endoscopist | -168
given oral antibiotics | -168
no improvement | -168
dysphonia | 0
cough | 0
deterioration of general condition | 0
body temperature 39 °C | 0
white blood cell count 18,900/mm3 | 0
hemoglobin level 11.3 g/dL | 0
CRP 64 ng/ml | 0
plasma glucose level 680 mg/dl | 0
pH 7.4 | 0
plasma osmolarity 320 mOsm/kg | 0
diagnosed as nonketotic hyperosmolar coma | 0
taken into intensive care unit | 0
intravenous insulin | 0
0.9 NaCl administered | 0
wide spectrum prophylactic antibiotic ceftriaxon 2 gr/day | 0
fever remained high | 72
neck ultrasound examination | 72
abscess formation in upper mediastinum | 72
cervicothoracic computed tomography (CT) | 72
gas and abscess formation in upper mediastinum | 72
pleural effusion in both hemithorax | 72
Gram stain of needle aspiration | 72
polymorphonuclear leukocytes existence | 72
no bacteria | 72
needle aspirate culture failed to show bacterial growth | 72
ceftriaxon discontinued | 72
meropenem 3 gr/day | 72
symptoms resolved | 120
control cervicothoracic CT | 240
abscess formation and pleural effusion almost disappeared | 240
discharged | 360