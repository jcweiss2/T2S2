53 years old | 0  
    male | 0  
    hypertension | 0  
    type 2 diabetes mellitus | 0  
    alcohol abuse | 0  
    massive bout of alcohol intake | -96  
    liquid diarrhoea | -96  
    self-medication by NSAIDs (ibuprofen) | -96  
    febrile respiratory distress | 0  
    diffuse cutaneous marbling | 0  
    emergency admission | 0  
    blood pressure preserved (mean blood pressure 70-80 mmHg) | 0  
    oxygen saturation 83% without oxygen therapy | 0  
    confused | 0  
    marbling involved all four members with purpuric lesions on the extremities | 0  
    oligo-anuric | 0  
    initiation of massive fluid infusion | 0  
    acute renal failure | 0  
    serum creatinine 4.7 mg/dL | 0  
    blood urea nitrogen 8.4 mmol/L | 0  
    severe inflammation | 0  
    C reactive protein 300 mg/L | 0  
    procalcitonin 195 mg/L | 0  
    metabolic acidosis (pH 7.24, bicarbonataemia 14 mmol/L) | 0  
    hyperlactataemia (6 mmol/L) | 0  
    liver enzymes TGO/TGP 1.5-2 N | 0  
    anemia (9.6 g/dL) | 0  
    subnormal platelet count (130 G/L) | 0  
    hyperleucocytosis (24 G/L) | 0  
    increased lactate dehydrogenase (800 UI/L) | 0  
    free bilirubin 25 mmol/L | 0  
    haptoglobinaemia normal 1.3 g/L | 0  
    schizocytosis 2% | 0  
    prothrombin time 15 s | 0  
    fibrinogen 6.1 g/L | 0  
    troponin 618 ng/mL | 0  
    chest X-ray showed pneumonia of the lower right lobe | 0  
    echocardiography demonstrated global left ventricle hypokinesia | 0  
    ejection fraction 20% | 0  
    probabilist antibiotherapy (ceftriaxone/levofloxacin) | 0  
    haemodialysis initiated | 0  
    severe pneumonia | 0  
    complicated by acute renal failure | 0  
    myocarditis | 0  
    pneumococcal infection confirmed by positive urinary pneumococcal antigenuria | 0  
    blood cultures negative | 0  
    after 2 days of supportive treatment and antibiotherapy | 48  
    still oligo-anuric | 48  
    confused | 48  
    cutaneous necrotic lesions appeared on extremities, legs, hands, thorax, nose | 48  
    skin biopsy in the necrotic zone showed fibrin thrombi and epidermolysis | 48  
    haemoglobinaemia dropped from 9.6 g/dL to 8.2 g/dL | 48  
    platelets dropped from 130 G/L to 60 G/L | 48  
    schizocytes rose to 4% | 48  
    haptoglobin decreased to <0.1 g/L | 48  
    situation worsened | 48  
    plasmatic exchanges (PE) initiated with plasma substitution | 96  
    after 4 days of PE | 168  
    renal function unchanged | 168  
    haemolysis parameters unchanged | 168  
    persistence of anuria | 168  
    haptoglobin <0.1 g/L | 168  
    severe thrombopenia (32 G/L) | 168  
    schizocytosis 11% | 168  
    skin lesions rapidly worsened with necrosis extension | 168  
    confusion persisted | 168  
    obnubilation persisted | 168  
    cardiac parameters improved | 168  
    troponin-ultrasensible decreased to 106 ng/mL | 168  
    improved left ventricular function (ejection fraction 30-35%) | 168  
    ECZ treatment initiated (first dose 1200 mg) | 168  
    ECZ 900 mg weekly for three doses | 168  
    three days after first ECZ injection | 216  
    mental confusion regressed | 216  
    rise in platelet count (48 G/L) | 216  
    haptoglobin plasma level 0.4 g/L | 216  
    platelets >150 G/L on day 6 | 216  
    diuresis resumed on day 10 | 240  
    renal function improved gradually | 240  
    dialysis withdrawal on day 14 | 336  
    renal function fully recovered (serum creatinine 0.8 mg/mL) | 600  
    ECZ therapy maintained at 1200 mg twice monthly | 600  
    skin lesions on nose and hands healed without sequelae | 600  
    legs and feet infected | 600  
    trans-tibial bilateral amputation necessary at 3 months | 2160  
    investigations into cause of TMA found normal ADAMTS13 activity | 2160  
    no monoclonal gammapathy | 2160  
    HIV negative | 2160  
    hepatitis C negative | 2160  
    Parvovirus B19 negative | 2160  
    cytomegalovirus serology negative | 2160  
    stool culture negative for STEC | 2160  
    PCR stools negative for shigatoxin genes | 2160  
    direct Coombs’ test positive | 2160  
    indirect Coombs’ test positive | 2160  
    plasma levels of complement factors normal | 2160  
    C3 824 mg/L | 2160  
    C4 119 mg/L | 2160  
    CH50 145% | 2160  
    normal activity of CAP regulators | 2160  
    CFI 106% | 2160  
    CFH 101% | 2160  
    CD46 leucocyte expression 13.6% | 2160  
    plasmatic C5b9 normal 63 ng/mL | 2160  
    screening for anti-CFH antibodies negative | 2160  
    genetic screening negative for complement gene variants | 2160  
    ECZ discontinued after 6 months | 4320  
    one year later | 8760  
    all biological parameters normal | 8760  
    serum creatinine 0.89 mg/dL | 8760  
    