25 years old | 0
female | 0
pregnant | 0
admitted to the hospital | 0
heart failure | 0
ventricular tachycardia | 0
complete atrioventricular canal repair | -7300
mitral regurgitation | -7300
left ventricular ejection fraction of 33% | -7300
mechanical mitral prosthesis implantation | -2190
cardiac resynchronization therapy | -2190
New York Heart Association Class III | -2190
unplanned pregnancy | -196
refused to terminate pregnancy | -196
carvedilol | -196
furosemide | -196
warfarin | -196
INR levels between 3.0 and 3.5 | -196
worsening heart failure | -84
hospitalization | 0
sore throat | 8
cough | 8
COVID-19 test result positive | 8
non-contrast chest computed tomography scan | 8
bilateral ground-glass opacities | 8
fever | 12
pulse oximetry oscillating between 89% and 93% SaO2 | 12
progressive reduction of arterial pressure | 12
foetal distress signs | 12
emergency caesarean delivery | 12
healthy premature baby | 12
negative RT-PCR test for SARS-CoV-2 infection | 12
progressive multisystem organ failure | 15
septic shock | 15
inflammatory and prothrombotic biomarkers | 15
severe impairment of the pulmonary parenchyma | 15
ventilation in volume control mode | 15
antibiotic therapy | 15
amiodarone | 15
methylprednisolone | 15
therapeutic unfractionated heparin | 15
inotropic drugs | 15
gradual clinical improvement | 30
extubated | 30
non-invasive support | 30
nasal oxygen catheter | 30
massive bleeding from the digestive tract and airways | 37
tachypnoea | 37
tachycardia | 37
respiratory failure | 37
re-intubation | 37
cardiopulmonary arrest | 37
death | 37
diffuse alveolar damage | 37
viral cytopathic effects | 37
small pulmonary thrombi | 37
acute tubular necrosis | 37
cerebral oedema | 37
villous maturation | 37
syncytial knots | 37
fibrin depositions | 37
central and peripheral acute placental infarcts | 37