54 years old | 0
    male | 0
    smoking | -40320
    hypothyroidism | -40320
    T2N2bM0 HPV+ SCC of left base of tongue | -40320
    metastases to cervical lymph nodes | -40320
    enrolled in OPTIMA trial | -40320
    received carboplatin/abraxane induction chemotherapy (cycle 1) | -40320
    complete resolution of primary tongue tumor | -40320
    decrease in size of cervical lymph nodes | -40320
    minimal side effects from chemotherapy | -40320
    admitted for inpatient chemoradiotherapy | 0
    received 5-FU | 0
    received paclitaxel | 0
    received hydroxyurea | 0
    developed fever | 0
    pancytopenia | 0
    intractable diarrhea | 0
    vomiting | 0
    pancytopenia refractory | 0
    hydroxyurea dose decreased | 0
    hydroxyurea held | 0
    clinical course worsened | 0
    developed septic shock | 0
    progressive desquamative skin lesions | 0
    acute kidney failure | 0
    sustained pancytopenia | 0
    persistent hemodynamic instability | 0
    requiring multiple vasopressors | 0
    hypoxia | 0
    transferred to ICU | 0
    intubated | 0
    transitioned to comfort care | 0
    expired | 288
    skin lesions involving head, chest, back, right arm | 288
    toxic epidermal necrolysis | 288
    bone marrow hypocellular (<5%) | 288
    diminished trilineage hematopoiesis | 288
    no megakaryocytes | 288
    diffuse acute tubular necrosis | 288
    gastrointestinal tract pale-appearing | 288
    severely damaged mucosa | 288
    Stenotrophomonas maltophilia positive cultures | 288
    DPYD*2A/c.1905+1G>A mutation | 288
    homozygosity confirmed | 288
