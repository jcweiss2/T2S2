79 years old | 0\
male | 0\
hypertension | -672\
ischemic heart disease | -672\
severe symptomatic aortic stenosis | -672\
aortic valve area 0.6 cm2 | -672\
transvalvular maximal and mean gradients 61 and 33 mm Hg | -672\
left ventricular ejection fraction of 45% | -672\
coronary artery bypass graft surgery | -5280\
mitral valve repair | -5280\
admitted to the hospital | 0\
transcarotid approach | 0\
TEE probe placed | 0\
SAPIEN 3 valve deployed | 0\
postprocedural TEE | 0\
prosthesis in good position | 0\
no visible paravalvular leak | 0\
gastric aspiration with an orogastric tube | 0\
blood-tinged secretions | 0\
extubated | 0\
transferred to the intensive care unit | 0\
chest pain | 2\
shivering | 2\
CT with intravenous contrast | 2\
pneumomediastinum | 2\
right hydropneumothorax | 2\
esophageal perforation suspected | 2\
right thoracic drain inserted | 2\
serosanguinous liquid drained | 2\
esophagogastroscopy | 2\
4-cm vertical perforation of the middle third of the esophagus | 2\
returned to the operating room | 7\
right thoracotomy | 7\
repair of an esophageal perforation | 7\
lysis of extensive pleural adhesions | 7\
esophageal laceration site found | 7\
large vertebral osteophyte visualized | 7\
primary closure of the esophageal wall | 7\
intercostal muscular flap mobilized | 7\
thoracic drains left in place | 7\
transferred to the intensive care unit | 7\
pneumonia | 24\
severe delirium | 24\
congestive heart failure | 24\
pulmonary edema | 24\
died | 720