4 years old | 0
male | 0
admitted to the emergency room | 0
fever | -72
abdominal pain | -72
neck pain | -72
trauma to the back of his skull | -96
grunting | 0
poor perfusion | 0
severe neck pain | 0
temperature 39 °C | 0
heart rate 200 per minute | 0
blood pressure 111/79 mmHg | 0
respiratory rate 40 per minute | 0
intravenous line inserted | 0
intravenous fluid administered | 0
septic work-up done | 0
broad spectrum antibiotics started | 0
admitted to the pediatric intensive care unit | 0
progressive left neck pain | 12
neck swelling | 12
lateral neck radiograph taken | 12
thickened prevertebral soft tissue | 12
computed tomography scan of the neck with contrast | 12
minimal fluid collection in the retropharyngeal space | 12
no definite abscess | 12
left jugular vein filling defect | 12
partial thrombosis of the left internal jugular vein | 12
brain venogram computed tomography | 12
thrombosis confirmed | 12
blood culture positive for Methicillin-sensitive Staphylococcus aureus (MSSA) | 24
repeated culture positive for MSSA | 48
cerebrospinal fluid culture negative | 24
echocardiography done | 48
no vegetation or signs of infective endocarditis | 48
diagnosis of Lemierre syndrome | 48
new left-sided neck swelling | 72
left vertebral artery aneurysm | 72
coiling of the aneurysm | 72
insertion of a peripherally inserted central catheter (PICC) line | 72
episodes of bradycardia | 72
ECG done | 72
Type I Brugada syndrome pattern | 72
elevated J point | 72
coved ST segment | 72
inverted T wave in precordial leads | 72
follow-up ECGs repeated | 96
abnormal ECG findings disappeared | 120
no family history of cardiac diseases or sudden death | 0
genetic studies for Brugada syndrome negative | 120
discharge from the hospital | 168
follow-up with pediatric cardiology | 168
counseled regarding the nature of Brugada syndrome | 168
ECGs repeated after discharge | 168
ECGs normal | 168
no findings of Brugada pattern | 168