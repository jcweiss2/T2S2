32 years old | 0
African American | 0
male | 0
admitted to the hospital | 0
bilateral lower extremities weakness | -48
inability to walk | -48
progressive bilateral lower extremities weakness | -2160
slurred speech | -336
deviation of the left eye | -336
hypothyroidism | -0
acquired immune deficiency syndrome | -0
CD4+ T-lymphocyte cell count <20 | -4320
plasma HIV RNA 206,000 | -4320
dysarthria | 0
horizontal nystagmus bilaterally | 0
dysmetria on finger-to-nose examination | 0
unsteady gait | 0
abnormal non-enhancing hyperintense T2 hypointense T1 signal | 0
lumbar puncture | 0
cerebrospinal fluid analysis | 0
hypoxic | 120
hypotensive | 120
altered mental status | 120
intubated | 120
broad-spectrum antibiotics | 120
transferred to the ICU | 120
VRE peri-rectal surveillance cultures | 120
negative VRE peri-rectal surveillance cultures | 120
failed multiple weaning attempts | 240
percutaneous tracheostomy | 240
percutaneous endoscopic gastrostomy tube placement | 240
severe watery diarrhea | 504
C. difficile glutamate dehydrogenase and toxin B tests | 504
positive C. difficile glutamate dehydrogenase and toxin B tests | 504
oral vancomycin | 504
diarrhea persisted | 672
bleeding per rectum | 672
digital rectal exam | 672
solid brown stool with specks old blood | 672
no fresh blood | 672
colonoscopy | 720
diffuse area of severely altered vascular, congested, erythematous, friable with contact bleeding | 720
hemorrhagic, inflamed, nodular, and ulcerated mucosa | 720
biopsies | 720
oral and rectal vancomycin with metronidazole | 720
blood culture | 720
no growth of any organism | 720
urine culture | 720
no growth of any organism | 720
tissue culture | 720
VRE | 720
echocardiogram | 720
no vegetation | 720
infectious disease consulted | 720
continue with oral and rectal vancomycin with metronidazole | 720
clinical condition improved | 840
diarrhea resolved | 840
discharged to a nursing home | 840