78 years old | 0
    male | 0
    admitted to the hospital | 0
    hydrocelectomy (Winkelmann's procedure) | -360
    scrotal pain | -360
    scrotal swelling | -360
    temperature of 38 degrees C | 0
    palpable peripheral pulses | 0
    leukocytosis (26000) | 0
    elevated CRP (300) | 0
    ultrasound revealed enlarged left testis | 0
    swelling and fluids in the scrotal content | 0
    enlarged epididymis | 0
    orchidoepididymitis | 0
    multiple abscesses | 0
    surgical exploration of the scrotum | 0
    left hemiscrotectomy | 0
    placement of suprapubic catheter | 0
    Actinomyces turicensis | 0
    Streptococcus viridans | 0
    Staphylococcus | 0
    necrosis | 0
    phlegmonous inflammation | 0
    abscesses of the scrotum | 0
    necrotizing fasciitis | 0
    hyperbaric oxygen chamber | 0
    parenteral administration of Imipenem 3 g daily | 0
    parenteral administration of Cefotaxim 6 g daily | 0
    parenteral administration of Metronidazol 2 g daily | 0
    intensive care unit management | 0
    resolution of critical condition | 0
    Mesh-Grafting | 0
    vacuum assisted closure | 0
    skin auto transplantation | 0
    