35 years old | 0
male | 0
height 169 cm | 0
weight 240 kg | 0
BMI 84 | 0
left leg pain | -24
redness | -24
swelling | -24
visited Department of Dermatology | -24
focused enhanced CT of left leg | -24
ruled out deep venous thrombosis | -24
cellulitis | -24
sent home | -24
prescription for Cefdinir | -24
symptoms deteriorated | -24
re-visited Department of Dermatology | -24
biochemistry analysis | -24
multiple organ dysfunction | -24
consulted our department | -24
history of recurrent cellulitis | -24
obese since childhood | -24
employed in home demolition | -24
unable to stand due to pain | 0
stretcher could not accommodate | 0
bed retrieved from ward | 0
nine people lifted onto bed | 0
side bars removed | 0
Glasgow Coma Scale score 15 | 0
blood pressure 174/65 mmHg | 0
heart rate 108 bpm | 0
respiratory rate 30 bpm | 0
SpO2 98% with 3 L/min oxygen | 0
body temperature 36.7℃ | 0
left leg redness | 0
left leg swelling | 0
tenderness | 0
venous gas analysis pH 7.352 | 0
PCO2 28.8 mmHg | 0
PO2 61.7 mmHg | 0
HCO3- 15.5 mmol/L | 0
lactate 6.2 mmol/L | 0
sinus tachycardia | 0
chest roentgenogram cardiac enlargement | 0
CT not performed due to equipment | 0
white blood cell count 6,800/μL | 0
neutrophil 96% | 0
lymphocyte 2% | 0
monocyte 2% | 0
hemoglobin 14.0 g/dL | 0
platelet count 9.0×104/μL | 0
C-reactive protein 12.8 mg/dL | 0
aspartate aminotransferase 315 IU/L | 0
alanine aminotransferase 93 IU/L | 0
glucose 78 mg/dL | 0
blood urea nitrogen 26.0 mg/dL | 0
creatinine 1.34 mg/dL | 0
creatinine phosphokinase 9,670 IU/L | 0
activated partial thromboplastin time 38.7 s | 0
international normalized ratio 1.83 | 0
fibrinogen 261 mg/dL | 0
fibrinogen degradation product 21.4 mg/dL | 0
tentative diagnosis of sepsis | 0
multiple organ failure | 0
left leg infection | 0
massive infusion of Ringer's lactate | 0
linezolid | 0
meropenem | 0
tracheal intubation | 0
surgical exploration of left leg | 0
necrotic soft tissue infection | 0
left leg amputation not performed | 0
nurses unable to reposition | 0
laboratory findings transiently improved | 24
oligouria continued | 0
cannula for renal replacement therapy impossible | 0
died of multiple organ failure | 96
culture of surgical material Streptococcus dysgalactiae | 0
blood culturing not performed | 0
super-super obesity | 0
