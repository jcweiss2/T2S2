64 years old | 0
woman | 0
right flank pain | -24
dysuria | -24
pollakuria | -24
non-contrast abdominopelvic CT revealed right renal pelvic stone | -24
diabetes | 0
hypertension | 0
hypothyroidism | 0
medications under control | 0
preoperative complete blood count | -24
preoperative serum urea | -24
preoperative creatinine | -24
preoperative ALT | -24
preoperative AST | -24
preoperative coagulation parameters | -24
preoperative urine culture | -24
underwent right PNL in prone position | 0
general anesthesia | 0
PNL started in lithotomy position | 0
ureteral catheter placement | 0
conversion to prone position |A0
collecting system visualized with contrast | 0
posterior middle calyx puncture between 11th and 12th ribs | 0
uncomplicated procedure | 0
16 Fr nephrostomy tube placement | 0
hemoglobin level 13 g/dl | 0
hemoglobin decreased to 11 g/dl | 0
respiratory distress during recovery | 24
referred to intensive care unit | 24
sudden severe hypotension | 24
900cc hemorrhagic fluid in drainage tube | 24
hemoglobin 8.1 g/dl | 24
postoperative tomography no hematoma | 24
postoperative tomography no adjacent organ injury | 24
nephrostomy tube clamped | 24
blood transfusion initiated | 24
two units erythrocyte suspension | 24
single unit fresh frozen plasma transfusion | 24
hemoglobin increased to 10 g/dl | 24
respiratory stabilization | 24
hemodynamic stabilization | 24
transferred to urology clinic | 24
serum aminotransferases rise end of first postoperative day | 24
LDH rise end of first postoperative day | 24
AST > 20 times ULN | 96
ALT > 25 times ULN | 96
LDH > 10 times ULN | 96
serum parameters normalized within 2 weeks | 336
discharged on postoperative 9th day | 216
ischemic hepatitis diagnosis established | 24
serum transaminases elevation 24 h after hypotension | 24
LDH elevation 24 h after hypotension | 24
normal serum bilirubin | 24
normal INR | 24
liver enzymes LDH decrease on 2nd day | 48
AST decrease on 6th day | 144
ALT decrease on 5th day | 120
normalization within 12th day | 288
hemorrhage after PNL | 24
intraoperative bleeding risk | 0
blood transfusion risk | 0
systemic hypotension secondary to hemorrhage | 24
hemorrhage contributed to ischemic hepatitis | 24
hypotension contributed to ischemic hepatitis | 24
routine serum biochemical parameters evaluation if hemorrhage suspected | 216
