Here is the table of events and timestamps:

65 years old | 0
female | 0
scheduled to undergo a left lobe hepatectomy | 0
hepatocelluar carcinoma | 0
liver cirrhosis | -672
chronic hepatitis B | -672
Child-Pugh class A | -672
premedication with glycoppyrolate | 0
general anesthesia induced with propofol, rocuronium, and remifentanil | 0
sevoflurane, remifentanil, and rocuronium for anesthesia maintenance | 0
intubated and ventilated mechanically | 0
monitored by EKG, arterial blood pressure, central venous pressure, and SpO2 | 0
stable vital signs | -1
sudden decrease in arterial blood pressure, end-tidal carbon dioxide, and SpO2 | -1
tachycardia and ST elevation on EKG | -1
diagnosed with VAE and PAE | -1
resuscitation with colloid and catecholamines | -1
massive air emboli in both left and right heart | -1
arterial blood gas analysis | -1
pH 7.278, pCO2 51.3 mmHg, PO2 84.6 mmHg, HCO3- 24.2 mmHg, SaO2 94.4% on FiO2 0.5 | -1
systolic blood pressure and heart rate maintained at approximately 90 mmHg and 110 beats/min | -10
central venous pressure approximately 2 mmHg | -10
end-tidal carbon dioxide restored to 32 mmHg | -10
arterial blood gas analysis | -30
pH 7.338, pCO2 44.3 mmHg, PO2 234.0 mmHg, HCO3- 24.0 mmHg, SaO2 99.6% on FiO2 1.0 | -30
norepinephrine infusion and fluid resuscitation | -30
air emboli in left heart disappeared | -100
hepatectomy restarted and completed | -100
systolic pressure maintained at approximately 90 mmHg | -100
total anesthesia time 5 hours | -100
2,950 ml of fluid administered | -100
total urinary output and blood loss 220 ml and 800 ml, respectively | -100
intubated and ventilated mechanically in ICU | -100
systolic pressure maintained at approximately 90 mmHg | -100
postoperative laboratory findings | -100
abnormal PT/PTT, fibrinogen, d-dimer, antithrombin III, CK-MB, and troponin-T | -100
postoperative EKG showed ST elevation in II, III, and aVF | -100
EKG findings recovered normally | -48
trans-thoracic echocardiogram showed unremarkable findings and no PFO | -48
vital signs stable | -48
norepinephrine infusion tapered out | -48
mental status unchanged | -240
brain CT and MRI revealed multiple acute cerebral infarctions | -240
weaned to Spontaneous ventilation with CPAP mode and extubated | -240
vital signs became unstable | -240
intravenous administration of catecholamines started | -240
panperitonitis confirmed by gram (+) cocci on peritoneal culture | -240
expired due to cardiac arrest caused by septic shock | -480