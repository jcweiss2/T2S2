27 years old | 0
female | 0
pregnant | 0
traveled to Southeast Asia | -8760
diarrhea | -448
abdominal pain | -336
watery diarrhea | -336
mucous bloody stools | -336
admitted to the hospital | 0
spontaneous preterm birth | 24
newborn died | 24
anemia | 0
hypoalbuminemia | 0
sigmoidoscopy | 0
reddish edematous mucosa | 0
mucopurulent exudate | 0
bacterial culture negative | 0
Clostridioides difficile toxin negative | 0
biopsy | 0
suspected severe ulcerative colitis | 0
transferred to hospital | 48
Glasgow Coma Scale score of E3V4M6 | 48
temperature of 37.3°C | 48
blood pressure of 150/100 mmHg | 48
pulse rate of 122 beats/min | 48
respiratory rate of 22 breaths/min | 48
percutaneous oxygen saturation of 92% | 48
distended abdomen | 48
peritoneal irritation | 48
anemia | 48
thrombocytopenia | 48
prolonged coagulation | 48
elevated inflammatory response | 48
hypoalbuminemia | 48
computed tomography | 48
edematous changes in the colorectum | 48
loss of haustra | 48
large amount of residue | 48
no megacolon | 48
no gastrointestinal perforation | 48
managed in ICU | 48
sigmoidoscopy | 48
pseudomembrane | 48
blood | 48
edematous mucosa | 48
faded reddish-purple mucosa | 48
biopsy | 48
emergency periodic acid-Schiff staining | 72
E. histolytica trophozoites | 72
diagnosed with fulminant amebic enteritis | 72
intravenous metronidazole | 72
ventilator management | 72
pulmonary edema | 72
inflammatory markers improved | 120
diarrhea disappeared | 120
fever disappeared | 120
weaned off ventilator | 120
diarrhea recurred | 480
fever recurred | 480
colonoscopy | 480
pseudomembrane disappeared | 480
punched-out ulcers | 480
CMV antigenemia test positive | 480
diagnosed with CMV enteritis | 480
intravenous ganciclovir | 480
symptoms improved | 504
laboratory data improved | 504
abdominal distension | 1440
colonoscopy | 1440
Gastrografin enema | 1440
severe stenosis | 1440
subtotal colectomy | 1440
ileorectal anastomosis | 1440
operative specimen | 1440
wall thickening | 1440
inflammation | 1440
stenosis | 1440
pathological examination | 1440
active inflammation | 1440
fibrosis | 1440
fibrotic stenosis | 1440
discharged | 4800