54 years old | 0
male | 0
Frontotemporal dementia (FTD) | 0
progressive abnormal emotional processing | 0
frontotemporal atrophy | 0
diagnosed with FTD | -87600
apathy | -87600
self-destructive impulsivity | -87600
weakness of lower limb | -87600
frequent syncope | -87600
fluctuation of blood pressure (BP) | -87600
taken anticholinergic drug | -87600
severe atrophy of bilateral frontal and temporal lobes | -87600
taken selective serotonin reuptake inhibitors | -87600
taken anticonvulsants | -87600
taken dopamine agonist | -87600
taken anticholinergic medications | -87600
anemia | 0
bleeding of stomach cancer | 0
hemoglobin 8.3 g/dl | 0
atrial fibrillation | 0
transferred to the operating room | 0
applied standard monitors | 0
BP 110/85 mmHg | 0
HR 85 beats/min | 0
administered thiopental 170 mg | 0
administered vecuronium 6 mg | 0
intubated successfully | 0
mechanical ventilation started | 0
tidal volume 450 ml | 0
respiration rate 10 breaths/min | 0
FIO2 0.5 | 0
end tidal CO2 30-35 mmHg | 0
anesthesia maintained with sevoflurane | 0
stable vital signs | 0
systolic/diastolic BP 110-130/708-90 mmHg | 0
HR 80-95 beats/min | 0
sudden drop in BP to 70/40 mmHg | 24
shedding 300 ml of blood | 24
atrial fibrillation at varying rates 110-130 beats/min | 24
administered 1500 ml Lactated Ringer's solution | 24
administered 1 unit packed red blood cells | 24
consulted cardiologist | 24
TEE performed | 24
TEE showed normal valves | 24
TEE showed contractility with adequate volume state | 24
no regional wall motion abnormality | 24
estimated ejection fraction 65% | 24
HR returned to 50 beats/min after synchronized cardioversion | 24
no change in BP | 24
bolus injection of ephedrine | 24
infused dopamine 10 µg/kg/min | 24
infused dobutamine 10 µg/kg/min | 24
infused norepinephrine 0.3 µg/kg/min | 24
no response to dopamine | 24
no response to dobutamine | 24
no response to norepinephrine | 24
high dose epinephrine 0.5-1.0 mg induced increasing BP | 24
used vasopressin 4 units/h after 10 units bolus dose | 24
BP returned to 110/65 mmHg | 24
HR returned to 75 beats/min | 24
infused dopamine 5 µg/kg/min | 24
infused dobutamine 5 µg/kg/min | 24
infused arginine vasopressin 4 U/h | 24
operation completed successfully | 24
transferred to intensive care unit | 24
titrated vasopressors | 24
stopped vasopressors completely at 24 h after surgery | 48
extubated | 48
transferred to general ward | 72
no sequelae | 72
