18 years old | 0
female | 0
8 weeks pregnant | 0
acute severe asthma | -720
short non-infective prodrome | -720
hypoxic cardiac arrest | -720
ventricular fibrillation | -720
resuscitation | -720
sinus tachycardia | -710
endotracheal intubation | -710
therapeutic hypothermia | -696
salbutamol | -696
ipratropium | -696
aminophylline | -696
hydrocortisone | -696
magnesium | -696
ketamine | -696
inhalation anesthesia with 1 MAC isoflurane | -696
severe hypercapnic acidosis | -696
neuromuscular blockade | -696
generalised status myoclonus | -48
ventilation improving | -48
intravenous sedatives ceased | -48
0.25–0.5 MAC isoflurane | -48
absent motor response to painful stimulus | 0
preserved pupillary reflexes | 0
preserved corneal reflexes | 0
preserved cough reflexes | 0
preserved gag reflexes | 0
spontaneously breathing | 0
severe generalised status myoclonus | 0
refractory to three antiepileptic medications | 0
electroencephalography | 0
generalised periodic discharges | 0
absent background rhythm | 0
reversible causes of coma eliminated | 0
biochemical causes eliminated | 0
metabolic causes eliminated | 0
septic causes eliminated | 0
drugs causes eliminated | 0
no shortness of breath | 0
denies chest pain | 0
no agreement about her neurological outcome | 8
additional social issues | 8
intensive social work support | 8
plasma neuron-specific enolase | 10
51 mcg/L | 10
somatosensory-evoked potential | 10
unhelpful due to myoclonus motion artefacts | 10
brain magnetic resonance imaging | 10
bilateral basal ganglia and frontoparietal cortex infarction | 10
extubated | 10
died in 24 h | 34