43 years old | 0
Hispanic female | 0
admitted to the hospital | 0
right upper quadrant abdominal pain | -168
fever | -168
nausea | -168
vomiting | -168
diarrhea | -168
hypotensive | 0
tachycardic | 0
temperature of 38.0 °C | 0
pulse of 138 beats per minute | 0
respiratory rate of 18 per minute | 0
blood pressure of 90/54 mm Hg | 0
pulse oximetry of 99% on room air | 0
dry mucosal membranes | 0
diffuse abdominal tenderness | 0
transferred to the intensive care unit | 0
septic shock | 0
white blood cell count of 5,620/µL | 0
hemoglobin of 11.7 g/dL | 0
sodium level of 130 mmol/L | 0
potassium of 3.3 mmol/L | 0
creatinine of 3.3 mg/dL | 0
glomerular filtration rate of 15.26 mL/min | 0
total bilirubin of 1.5 mg/dL | 0
aspartate aminotransferase of 246 U/L | 0
alanine aminotransferase of 185 U/L | 0
alkaline phosphatase of 131 U/L | 0
lipase of 35 U/L | 0
lactic acid of 7.2 mmol/L | 0
COVID-19 positive | 0
CT scan of the abdomen | 0
poorly defined hypodense cystic structure in the right liver lobe | 0
ultrasound | 0
9.9-cm mass in the right lobe of the liver | 0
MRI scan of the abdomen | 0
heavily septated 13-cm hepatic abscess in the posterior right hepatic lobe | 0
intravenous vancomycin | 0
piperacillin/tazobactam | 0
percutaneous drainage | 0
1,110 mL of purulent fluid | 0
Streptococcus viridans | 0
switched to ampicillin/sulbactam | 0
RUQ pain improved | 0
discharged | 192
left lower quadrant abdominal pain | 192
repeat CT of the abdomen | 192
decreased size of the liver lesion | 192
pelvic abscess measuring 13.6 × 5 cm | 192
unchanged pneumoperitoneum | 192
perforated sigmoid diverticulum | 192
CT-guided percutaneous drainage | 192
mixed gram-positive and gram-negative flora | 192
Candida albicans | 192
amoxicillin | 192
fluconazole | 192
drain removal | 240
improvement of LLQ pain | 240