38 years old | 0
female | 0
13th week of pregnancy | 0
abdominal discomfort | -24
nausea | -24
vomiting | -24
no fever | -24
no vaginal discharge | -24
admitted to the ER | 0
discharged home | 0
persistent abdominal pain | 144
nausea | 144
vomiting | 144
tachycardic | 144
diffuse abdominal pain | 144
guarding on the right quadrants | 144
neutrophilia | 144
low prothrombinemia | 144
acute renal failure | 144
high procalcitonin | 144
high c-reactive protein | 144
moderate fluid in all quadrants | 144
good foetal vitality | 144
hypotension | 144
general abdominal guarding | 144
hyperlacticaemia | 144
hypokalaemia | 144
hyperglycaemia | 144
septic shock | 144
emergency exploratory laparotomy | 144
generalised purulent peritonitis | 144
perforated acute appendicitis | 144
appendicectomy | 144
abdominal washing | 144
laparostomy | 144
admitted to the ICU | 144
septic shock | 144
need for vasopressor therapy | 144
need for dialysis | 144
intravenous piperacillin-tazobactam | 144
laparostomy revision | 192
marked bowel oedema | 192
bowel distention | 192
mild intraabdominal soiling | 192
peritoneal lavage | 192
new laparostomy | 192
progressive closure technique | 192
surgical revision | 216
abdominal cavity primary closed | 216
antibiotherapy adjusted | 216
piperacillin-tazobactam suspended | 216
amoxicillin with clavulanic acid | 216
transferred to the obstetrics ward | 288
discharged home | 336
elective caesarean section | 1008
gave birth to a healthy child | 1008
ventral hernia | 1092