54 years old | 0  
    female | 0  
    type 2 diabetes mellitus | 0  
    end-stage renal disease | 0  
    presented to the emergency department | 0  
    headache | -240  
    photophobia | -240  
    chronic cough | -240  
    weight loss | -240  
    low-grade fever | -240  
    close contact with tuberculosis | -26160  
    febrile | 0  
    tachycardic | 0  
    mild impairment of alertness | 0  
    diffuse crackles | 0  
    left lung | 0  
    white blood cell count 4800 cells/μL | 0  
    absolute lymphocyte count 816 cells/μL | 0  
    hemoglobin 10.3 g/dL | 0  
    blood sugar 111 mg/dL | 0  
    normal liver function tests | 0  
    creatinine 7.2 mg/dL | 0  
    blood urea nitrogen 59 mg/dL | 0  
    bilateral interstitial infiltrates | 0  
    multiple ring-shaped lesions | 0  
    posterior areas of both hemispheres | 0  
    acid-fast bacilli sputum culture positive | 0  
    Mycobacterium tuberculosis complex | 0  
    no antibacterial resistance | 0  
    HIV1/2 negative | 0  
    toxoplasma serologies negative | 0  
    opening pressure 30 cm H2O | 0  
    red blood cell count 1000 cells/μL | 0  
    WBC 114 cells/μL | 0  
    lymphocytes 92% | 0  
    glucose 30 mg/dL | 0  
    proteins 161 mg/dL | 0  
    CSF neurocysticercosis serology negative | 0  
    cryptococcal antigen negative | 0  
    CSF Mycobacterium tuberculosis stain negative | 0  
    CSF culture negative | 0  
    adenosine deaminase negative | 0  
    PCR positive for MTB | 0  
    anti-TB therapy started | 0  
    rifampin | 0  
    isoniazid | 0  
    pyrazinamide | 0  
    ethambutol | 0  
    pyridoxine | 0  
    adjunctive dexamethasone | 0  
    mental status deteriorated | 24  
    admission to intensive care unit | 24  
    initiation of hemodialysis | 24  
    uremia | 24  
    clinical improvement | 24  
    acute abdominal pain | 504  
    hematemesis | 504  
    CT abdomen loculated multiseptated gas | 504  
    fluid collection gastric fundus | 504  
    free intra-abdominal air | 504  
    gastric perforation | 504  
    exploratory laparotomy | 504  
    complete stomach necrosis | 504  
    total gastrectomy | 504  
    intestinal discontinuity | 504  
    cervical esophagostomy | 504  
    jejunostomy tube placement | 504  
    oral anti-TB switched to intravenous | 504  
    amikacin | 504  
    linezolid | 504  
    levofloxacin | 504  
    rifampin continued | 504  
    septic shock | 504  
    intubation | 504  
    mechanical ventilation | 504  
    empiric piperacillin-tazobactam | 504  
    vascular thrombosis | 504  
    broad irregularly branched hyphae | 504  
    angio-invasive gastric mucormycosis | 504  
    acid-fast bacilli stain negative | 504  
    culture negative | 504  
    liposomal amphotericin B initiated | 504  
    TB treatment maintained | 504  
    isoniazid plus rifampin continued | 672  
    liposomal amphotericin B switched to posaconazole | 672  
    clinical stabilization | 672  
    improvement | 672  
    returned to Latin America | 672  
    gastrointestinal mucormycosis | 0  
    disseminated tuberculosis | 0  

