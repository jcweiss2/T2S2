47 years old | 0
    obese | 0
    short neck | 0
    body mass index 42 kg/m2 | 0
    admitted in ED | 0
    respiratory distress | 0
    asphyxiation | 0
    twenty-sixth postoperative day after total thyroidectomy | 624
    history of present illness | -624
    total thyroidectomy | -624
    fine-needle biopsy confirmed medullary thyroid carcinoma | -624
    enlarged fibrotic multinodular massive goiter | -624
    tracheal compression | -624
    preoperative neck stiffness | -624
    preoperative throat fullness | -624
    preoperative hoarseness | -624
    preoperative orthopnea | -624
    preoperative difficulty breathing | -624
    transferred to post anesthesia care unit | -624
    tracheostomy tube in place | -624
    extensive neck dissection | -624
    difficult neck dissection | -624
    presumed RLN injury | -624
    intraoperative tracheomalacia | -624
    postoperative period unremarkable | -624
    discharged from hospital | -624
    second postoperative day | 48
    next six days | 168
    gradual neck stiffness | 168
    gradual throat tightness | 168
    gradual dyspnea | 168
    pain during swallowing | 168
    subfebrile condition | 168
    cough | 168
    purulent sputum | 168
    existing tracheostomy | 168
    suspected tracheostomy tube problem | 168
    referred to otorhinolaryngologist | 168
    indirect mirror laryngoscopy | 168
    right VCP | 168
    neck visibly swollen | 168
    reddish neck color | 168
    new onset dyspnea | 168
    postoperative course not considered | 168
    possibility of surgical complications not considered | 168
    decannulate | 168
    discharge patient | 168
    continued worsening of complaints | 168
    breathing difficulties worsening | 168
    referred to pulmonologist | 168
    increased bronchodilators dosages | 168
    no clinical improvement | 168
    hypertension | -8760
    COPD | -8760
    regular Indapamide | -8760
    regular Candesartan | -8760
    regular Albuterol | -8760
    regular Tiotropium bromide | -8760
    critical condition | 0
    tripod position | 0
    severe tachy-dyspnea | 0
    respiratory rate 48/min | 0
    desaturation SpO2 68% | 0
    intense cyanosis | 0
    orthodeoxia | 0
    orthopnea | 0
    biphasic stridor | 0
    increased work of breathing | 0
    diaphoresis | 0
    impossible swallowing | 0
    tachycardia 144 beats/min | 0
    hypertension 186/110 mmHg | 0
    aphonia | 0
    temperature 38.9 ℃ | 0
    post thyroidectomy scar reddish | 0
    tracheostomy obliterated | 0
    large submandibular mass | 0
    painful submandibular mass | 0
    bilateral expiratory rhonchi | 0
    purulent sputum | 0
    reddish skin discoloration | 0
    contrast enhanced CT scan of neck | 0
    large pre-tracheal cavity | 0
    spongiform appearance | 0
    gaseous content | 0
    closed glottis | 0
    immobile glottic musculature | 0
    bilateral VCP | 0
    cannot intubate cannot ventilate scenario | 0
    pre-oxygenation with 100% O2 | 0
    SpO2 78% | 0
    rapid sequence induction | 0
    fentanyl 200 µg | 0
    propofol 300 mg | 0
    succinylcholine 100 mg | 0
    Cormack Lehane 2a grade | 0
    closed vocal cords | 0
    small cleft posteriorly | 0
    endotracheal tube 5.5 ID | 0
    uneventful ventilation | 0
    re-tracheostomy | 0
    pre-tracheal fascia opened | 0
    stench of decay | 0
    gossypiboma | 0
    abscess cavity cultures Streptococcus viridans | 0
    ARDS ruled out | 0
    preserved lung parenchyma | 0
    extensive antimicrobial course | 0
    cured | 0
    discharged | 24
    decannulated after a month | 720
    full recovery from neck inflammation | 720
    gradual voice rehabilitation | 720
    voice fatigue | 2928
    ethical approval | -624
    written informed consent | -624
    CREC 2022/166 approval | -624
    