57 years old | 0
female | 0
chronic congestive heart failure | -8760
postpartum cardiomyopathy | -8760
type 2 diabetes | -8760
hypothyroidism | -8760
admitted to the hospital | 0
acute respiratory failure | 0
cardiogenic shock | 0
new-onset nonischemic cardiomyopathy | 0
left ventricular ejection fraction (LVEF) drop | 0
worsening preexisting hypokalemia | 0
loop diuretics | 0
spironolactone | 0
losartan | 0
elevated serum morning cortisol | 0
elevated ACTH | 0
low aldosterone/renin ratio | 0
high 24-hour free urine cortisol | 0
DHEA sulfate levels | 0
Metanephrine plasma levels | 0
CT abdomen | 0
symmetrical enlargement of both adrenal glands | 0
endocrinology consultation | 0
denies recent weight gain | 0
denies headaches | 0
denies vision change | 0
denies abdominal striae | 0
denies proximal muscle weakness | 0
denies hirsutism | 0
denies acne | 0
denies history of kidney stones | 0
denies steroid use | 0
normal blood pressure | 0
no cushingoid features | 0
normal pituitary gland | 0
stress-induced cardiomyopathy | 0
vasopressors | 0
diuretics | 0
improved cardiac condition | 168
near resolution of adrenal enlargement | 168
normalization of morning cortisol | 168
normalization of ACTH levels | 168
normalization of 24-h free urine cortisol | 168
normalized potassium levels | 168
improvement in LVEF | 168
discharged from the hospital | 168
lost to endocrinology follow-up | 720
cortisol and ACTH checks within normal limits | 1008
readmitted to the hospital | 2160
septic shock | 2160
pneumonia | 2160
worsening cardiac failure | 2160
liver failure | 2160
gastrointestinal bleeding | 2160
died | 2160
normal morning cortisol level | 2160
no autopsy | 2160
dobutamine | 0
milrinone | 0
diuresis with IV bumetamide | 0
transitioned to oral bumetamide | 24