74 years old | 0\
male | 0\
hypertension | 0\
diabetes mellitus | 0\
intermittent subjective fever | -96\
rigors | -96\
generalized headache | -96\
altered mentation | -96\
body malaise | -96\
nausea | -96\
vomiting | -96\
febrile | 0\
tachypneic | 0\
disoriented | 0\
tachycardic | 0\
low blood pressure | 0\
saturating at 98% on room air | 0\
normal vesicular breath sounds | 0\
normal abdominal examination | 0\
intravenous (IV) resuscitation | 0\
analgesia | 0\
white blood cell count (WBC) of 8.2 × 103/μL | 0\
hemoglobin (Hb) of 11.5 g/dL | 0\
thrombocytopenia of 46,000/mm3 | 0\
elevated creatinine 117 μmol/L | 0\
BUN 10.5 mmol/L | 0\
low sodium of 131 mmol/L | 0\
normal serum electrolytes | 0\
normal liver | 0\
normal coagulation profile | 0\
normal Chest X-ray | 0\
P. falciparum with high parasitemia | 0\
admitted to the intensive care unit (ICU) | 0\
intravenous artesunate-based regimen | 0\
supportive measures | 0\
shifted to the general ward | 72\
acute abdomen | 120\
progressive, dull, constant generalized abdominal pain | 120\
nausea | 120\
non-bilious vomiting | 120\
anxious | 120\
afebrile | 120\
diaphoretic | 120\
tachycardic | 120\
tachypneic | 120\
hypotensive | 120\
saturating well on room air | 120\
distended abdomen | 120\
tender on superficial palpation | 120\
inaudible bowel sounds | 120\
low Hb of 7.1 g/dL | 120\
hypoechoic nodular cystic area | 120\
hyperdense intrasplenic hematoma | 120\
hypodense subcapsular hematoma | 120\
splenic laceration | 120\
intraperitoneal free fluid | 120\
grade 3 splenic injury | 120\
blood products | 120\
adequate resuscitation | 120\
explorative laparotomy | 120\
splenectomy | 120\
2.5 L of frank blood | 120\
enlarged spleen | 120\
long laceration on the upper pole | 120\
uneventful postoperative period | 168\
discharged home | 168