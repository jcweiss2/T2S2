37 years old|0
female|0
admitted to the hospital|0
poorly controlled type 2 diabetes mellitus|0
peripheral neuropathy|0
morbid obesity|0
BMI of 45.8 kg/m2|0
obstructive sleep apnea|0
gastroesophageal reflux disease|0
depression|0
intellectual disability|0
metformin 500 mg twice a day|0
hemoglobin A1c was 9.8%|0
sitagliptin added|0
canagliflozin added|0
pain in the left gluteal region|-672
dysuria|-672
trimethoprim/sulfamethoxazole initiated|-672
urinary tract infection|-672
urine culture not collected|-672
no improvement|-672
go to the hospital|-168
afebrile (36.9°C)|0
tachycardic (117 beats/minute)|0
blood pressure of 144/79 mmHg|0
respiratory rate of 19 breaths/minute|0
lethargic|0
distress|0
suprapubic tenderness|0
induration to the left gluteal region|0
perineum induration|0
blood glucose of 402 mg/dL|0
serum bicarbonate of 12 mmol/L|0
elevated anion gap of 24 mmol/L|0
lactate of 1.8 mmol/L|0
serum electrolytes within normal range|0
creatinine within normal range|0
blood urea nitrogen within normal range|0
serum osmolarity of 295 mOsm/kg|0
glycosuria|0
ketonuria|0
glucose 4+|0
ketones 1+|0
b-hydroxybutyrate of 2.49 mmol/L|0
pH of 7.23|0
PCO2 of 34 mmHg|0
computed tomography of abdomen and pelvis|0
subcutaneous edema|0
air within medial left gluteal soft tissues|0
locules of air extending into presacral soft tissues|0
Fournier’s gangrene|0
intravenous normal saline 0.9% bolus|0
IV ceftazidime 2 g|0
IV clindamycin 600 mg|0
vancomycin 2 g|0
debridement|0
incision and drainage of left gluteal region|0
hypotensive|48
tachycardic|48
ongoing infection|48
sepsis|48
second surgical exploration|48
fluid resuscitation|48
admitted to surgical ICU|48
intubated|48
vasopressors required|48
antibiotics switched to vancomycin|48
piperacillin/tazobactam|48
surgical re-explorations|72
further debridement|72
laparoscopic transverse loop colostomy|168
fecal diversion|168
prevent further infection of perineum|168
DKA management|72
subcutaneous insulin|72
serum ketones identified|72
anion gap persisted|72
insulin infusion started|96
aggressive fluid resuscitation started|96
anion gap closed|120
acidosis resolved|120
transferred to general medical floor|408
discharged|672
urinary catheter|672
vacuum dressing|672
colostomy|672
short-term rehabilitation facility|672
insulin glargine 18 U started|672
discontinue canagliflozin|672
discontinue sitagliptin-metformin|672
