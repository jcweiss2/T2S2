33 years old | 0
female | 0
cachectic | 0
admitted to the hospital | 0
past medical history of untreated hepatitis C infection | -672
intravenous drug abuse | -672
acute respiratory failure | 0
mechanical ventilation | 0
MSSA bacteremia | 0
tricuspid valve endocarditis | 0
spontaneous right sided PTX | -240
chest tube placement | -240
temperature of 100.9 F | 0
pulse of 113/min | 0
respiratory rate of 18/min | 0
blood pressure of 109/65 mmHg | 0
pulse oximetry of 100% on FiO2 of 40% | 0
coarse breath sounds bilaterally in anterior lung fields | 0
3/6 systolic murmur best heard in the right lower sternal border | 0
chest tube in place | 0
resolution of PTX | 0
hemoglobin of 8.2 gm/dL | 0
white blood cell count of 10,000/mL | 0
platelet count of 52,000/mm3 | 0
BUN of 21 mg/dL | 0
creatinine of 0.48 mg/dL | 0
sodium of 138 mEq/L | 0
potassium of 3.6 mEq/L | 0
normal coagulation parameters | 0
persistent MSSA bacteremia | 0
pleural fluid cultures did not isolate any organism | 0
large, mobile, prolapsing 3.5 × 1.5 cm2 vegetation on the anterior leaflet of TV | 0
moderate tricuspid regurgitation | 0
bilateral septic emboli to lungs | 0
cavitary lesions | 0
small bilateral pleural effusions | 0
bibasilar infiltrates | 0
empiric antibiotics | 0
cardiothoracic surgery consultation | 0
septic shock | 24
acute renal failure | 24
urinary tract infection | 24
sudden onset respiratory distress | 240
new right sided PTX | 240
second chest tube placement | 240
not a suitable candidate for valve surgery | 240
recurrent noniatrogenic pneumothoraces | 240
three chest tubes on the right | 240
two chest tubes on the left | 240
comfort care measures | 336
died post terminal extubation | 336
autopsy not performed | 336