72 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
high-grade fever | -96 | 0 | Factual
influenza B virus infection | -96 | 0 | Factual
wife diagnosed with influenza B virus infection | -120 | -96 | Factual
daughters diagnosed with influenza B virus infection | -120 | -96 | Factual
rapid test positive for influenza B antigens | -96 | -96 | Factual
oseltamivir administered | -96 | -96 | Factual
persistent fever | -48 | 0 | Factual
dyspnea at rest | -48 | 0 | Factual
admitted to hospital | 0 | 0 | Factual
temperature 38.7°C | 0 | 0 | Factual
blood pressure 117/80 mmHg | 0 | 0 | Factual
heart rate 76 beats/min | 0 | 0 | Factual
oxygen saturation level 88% | 0 | 0 | Factual
fine crackles in lung fields | 0 | 0 | Factual
white blood cell count 7400/mm3 | 0 | 0 | Factual
C-reactive protein 18.1 mg/dL | 0 | 0 | Factual
aspartate transaminase 91 IU/L | 0 | 0 | Factual
L-lactate dehydrogenase 362 IU/L | 0 | 0 | Factual
creatine kinase 793 IU/L | 0 | 0 | Factual
Krebs von den Lungen-6 1772 U/mL | 0 | 0 | Factual
hypoxemia | 0 | 0 | Factual
arterial blood gas analysis | 0 | 0 | Factual
ground-glass opacity in lung fields | 0 | 0 | Factual
chest computed tomography | 0 | 0 | Factual
diffuse ground-glass opacity in lung fields | 0 | 0 | Factual
high-flow nasal oxygen support | 0 | 129 | Factual
intravenous peramivir | 0 | 129 | Factual
antibiotics | 0 | 129 | Factual
piperacillin/tazobactam | 0 | 129 | Factual
levofloxacin | 0 | 129 | Factual
reticular shadow on chest CT worsened | 72 | 72 | Factual
PaO2/FiO2 ratio deteriorated | 72 | 72 | Factual
severe ARDS | 72 | 129 | Factual
mechanical ventilation proposed | 72 | 72 | Factual
high levels of positive end-expiratory pressure proposed | 72 | 72 | Factual
patient refused intubation | 72 | 72 | Factual
polymyxin B-immobilized fiber column hemoperfusion | 72 | 72 | Factual
intravenous methylprednisolone | 144 | 144 | Factual
noninvasive positive pressure ventilation support | 144 | 129 | Factual
immunosuppressant therapy | 144 | 129 | Factual
intravenous cyclophosphamide | 144 | 129 | Factual
patient's condition worsened | 144 | 129 | Factual
patient died | 129 | 129 | Factual
autopsy performed | 129 | 129 | Factual
diffuse alveolar damage | 129 | 129 | Factual
prominent hyaline membranes | 129 | 129 | Factual
no specific abnormality in other organs | 129 | 129 | Factual
bacterial infection | 0 | 0 | Negated
fungal infection | 0 | 0 | Negated