56 years old | 0
male | 0
type 2 diabetes mellitus | 0
chronic obstructive pulmonary disease | 0
obstructive sleep apnea | 0
coronary artery disease | 0
heart failure with preserved ejection fraction | 0
tobacco abuse disorder | 0
alcohol use disorder | 0
presented to tertiary center critical care unit | 0
septic shock | 0
left lower extremity osteomyelitis | 0
found unresponsive | 0
intubated | 0
significant other found in apartment | 0
drinks 5 beers daily on weekdays | 0
increased alcohol use over last 3 months | -2160
eats frozen meals for last 3 months | -2160
blood cultures positive for methicillin-sensitive Staphylococcus aureus | 0
treated with appropriate antibiotics | 0
vascular surgery consulted | 0
no surgical intervention | 0
infectious diseases consulted | 0
admitted to ICU | 0
managed with pressor support | 0
managed with antibiotic treatment | 0
peculiar rash on presentation | 0
petechiae | 0
palpable hemorrhagic lesions | 0
rash resembling vasculitis | 0
rash on dorsal surfaces of hands | 0
rash on plantar surfaces of feet | 0
rash on legs | 0
rash on lips | 0
rash on gingiva | 0
rash present prior to antibiotics | 0
rash unchanged with antibiotics | 0
CBC normal white blood cell count | 0
hemoglobin slightly low | 0
MCV near normal | 0
platelet count within normal | 0
creatinine elevated | 0
coagulation factors normal | 0
ESR elevated | 0
C-reactive protein elevated | 0
immunologic workup pursued | 0
ANA negative | 0
ANCA IgG <1:20 | 0
Complement C3 elevated | 0
Complement C4 normal | 0
HIV negative | 0
hepatitis panel negative | 0
immunologic workup unremarkable | 0
nutritional deficiency considered | 0
plasma vitamin C levels drawn | 0
started on IV vitamin C | 0
vitamin C levels low | 0
diagnosed with scurvy | 0
skin findings improved | 168
mentation improved | 168
sepsis treatment | 0
inflammatory markers resolved | 168
creatinine resolved | 168
elevated ESR | 0
elevated C-reactive protein | 0
petechiae on plantar feet | 0
palpable lesions on dorsum of hands | 0
hyperkeratosis | 0
perifollicular hemorrhage | 0
gingival hemorrhage | 0
corkscrew hairs | 0
joint pain | 0
myalgias | 0
dry skin | 0
vasomotor instability | 0
vitamin C deficiency | 0
vitamin C treatment | 0
tube feeds started | 0
no ethical approval required | 0
informed consent obtained | 0
