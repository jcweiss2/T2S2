32 years old | 0
woman | 0
diagnosed with JAK2 mutation-negative essential thrombocythemia (ET) | -144000
treated by pipobroman for 7 years | -144000
treated by hydroxyurea for 4 years | -144000
treated by anagrelide for 3 years | -144000
began complaining about asthenia | -1464
gradual decrease in hemoglobin level | -1464
anagrelide stopped | -1464
bone marrow biopsy performed | -720
occurrence of grade 2 myelofibrosis | -720
hematologic tests revealed more than 20% blastic cells in peripheral blood | -504
ET with myelofibrosis evolved into acute myeloid leukemia | -504
received allogeneic bone marrow hematopoietic stem-cell transplantation (HSCT) | 0
admitted to intensive care unit (ICU) for acute respiratory distress syndrome (RDS) | 0
blood cultures yielded Staphylococcus aureus | 0
blood cultures yielded Escherichia coli | 0
broad-spectrum antibiotherapy (tazobactam/piperacillin, amikacin, vancomycin) | 0
furosemide for acute pulmonary edema | 0
rapid improvement of patient condition | 0
oral fluconazole prophylaxis (400 mg/day) started | 0
readmitted to ICU for acute RDS | 12
septic shock with no microbiological evidence of infection | 12
became afebrile after empirical antibiotherapy (ceftazidime, linezolid) | 12
presented with first symptoms of Graft-versus-Host Disease (GvHD) | 37
GvHD developed to skin | 37
GvHD developed to gastrointestinal tract | 37
GvHD developed to liver | 37
received corticosteroids | 37
received inolimomab | 37
received sirolimus | 37
received basiliximab | 37
digestive disorders remained chronic | 37
hemorrhagic manifestations | 37
readmitted to ICU for similar respiratory symptomatology | 63
new antibiotic regimen (imipenem, ciprofloxacin, ceftriaxone) | 63
intravenous caspofungin (50 mg/day) started | 63
routine microbiological surveillance cultures performed weekly | 63
Candida albicans isolated from oropharynx swab | -1464
Candida albicans isolated from rectal swab or stools | -1464
Candida albicans isolated from urine | -1464
Candida albicans no longer isolated | 0
colonization of gastrointestinal tract by C. kefyr | 0
colonization of urinary tract by C. kefyr | 0
increasing fungal load | 0
caspofungin stopped | 0
oral fluconazole (400 mg/day) restarted | 0
neutropenic patient suffered from unexplained fever | 0
thoracic computed tomography (CT) performed | 0
CT imaging showed pulmonary nodules suspected to be pulmonary aspergillosis | 0
antifungal therapy switched to voriconazole | 0
serum galactomannan (GM) assay performed twice a week | 0
GM assay index on bronchoalveolar lavage (BAL) was negative | 0
BAL culture yielded no Aspergillus | 0
BAL culture yielded heavy growth of C. kefyr | 0
blood cultures remained negative | 0
no other pathogen found | 0
measurement of (1→3)-β-d-glucan antigenemia revealed elevated serum concentration (411 pg/mL) | 0
possible deep candidiasis suspected | 0
treatment with caspofungin resumed | 0
follow-up CT showed increase in size and number of pulmonary lesions | 0
readmitted to ICU with acute renal failure | 0
died of multiple organ failure | 168
