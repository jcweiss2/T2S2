42 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
presented to the infectious diseases clinic | 0 | 0 | Factual
generalized weakness | -2160 | 0 | Factual
fever | -2160 | 0 | Factual
cough | -2160 | 0 | Factual
weight loss | -2160 | 0 | Factual
lived in Guatemala | -8760 | -2160 | Factual
sought medical attention in Guatemala | -2160 | -2160 | Factual
HIV-antibody test positive | -2160 | -2160 | Factual
sputum AFB smear positive | -2160 | -2160 | Factual
HIV-1 Western blot test positive | -168 | -168 | Factual
CD4 cell count 10/µL | -168 | -168 | Factual
HIV RNA titer 18,000 copies/mL | -168 | -168 | Factual
anti-tuberculosis medications started | -168 | -128 | Factual
isoniazid | -168 | -128 | Factual
rifampin | -168 | -128 | Factual
ethambutol | -168 | -128 | Factual
pyrazinamide | -168 | -128 | Factual
fluconazole | -168 | -128 | Factual
trimethoprim/sulfamethoxazole | -168 | -128 | Factual
generalized weakness persisted | -128 | 0 | Factual
fever persisted | -128 | 0 | Factual
admitted to KU hospital | 0 | 0 | Factual
body temperature 37.6℃ | 0 | 0 | Factual
oral thrush | 0 | 0 | Factual
hepatosplenomegaly | 0 | 0 | Factual
ascites | 0 | 0 | Factual
hemoglobin 10.6g/dL | 0 | 0 | Factual
white blood cell 2,700/µL | 0 | 0 | Factual
platelet 58,000/µL | 0 | 0 | Factual
total bilirubin 2.4mg/dL | 0 | 0 | Factual
AST/ALT 131/48IU/L | 0 | 0 | Factual
ALP 114IU/L | 0 | 0 | Factual
GGT 133 IU/L | 0 | 0 | Factual
chest X-ray showed costophrenic angle blunting | 0 | 0 | Factual
fluid shifting in the right hemithorax | 0 | 0 | Factual
mild pneumonic infiltration in left lung | 0 | 0 | Factual
disseminated tuberculosis suspected | 0 | 0 | Factual
Mycobacterium tuberculosis identified | 0 | 0 | Factual
anti-tuberculosis medication continued | 0 | 240 | Factual
anti-retroviral agents started | 0 | 0 | Factual
zidovudine | 0 | 120 | Factual
lamivudine | 0 | 120 | Factual
efavirenz | 0 | 120 | Factual
pancytopenia progressed | 24 | 120 | Factual
hemoglobin 7.4g/dL | 120 | 120 | Factual
white blood cell 1,070/µL | 120 | 120 | Factual
platelet 13,000/µL | 120 | 120 | Factual
rifampin discontinued | 120 | 120 | Factual
zidovudine discontinued | 120 | 120 | Factual
trimethoprim/sulfamethoxazole discontinued | 120 | 120 | Factual
new pulmonary infiltrates | 120 | 120 | Factual
septic shock | 120 | 120 | Factual
empirical antibiotic therapy started | 120 | 120 | Factual
piperacillin/tazobactam | 120 | 240 | Factual
transferred to intensive care unit | 144 | 144 | Factual
mechanical ventilator support | 144 | 240 | Factual
Gram stain and ordinary culture showed no pathologic organisms | 144 | 240 | Factual
bone marrow aspiration and biopsy performed | 216 | 216 | Factual
died | 240 | 240 | Factual
refractory septic shock | 240 | 240 | Factual
hypoxia | 240 | 240 | Factual
Histoplasma capsulatum identified | 240 | 240 | Factual
disseminated histoplasmosis confirmed | 240 | 240 | Factual