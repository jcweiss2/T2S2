54 years old | 0
male | 0
admitted to the hospital | 0
chronic cough | -672
squamous cell carcinoma | -672
ostium secundum atrial septal defect | -672
gastroesophageal reflux disease | -672
lung lobectomy | 0
general anesthesia | 0
SpO2 96%-100% | 0
left radial arterial and central venous pressures monitored | 0
video-assisted thoracoscopy | 0
left lower lobar pulmonary artery and inferior pulmonary vein division mobilized and stapled | 0
open thoracotomy | 0
seventh subcarinal lymph node dissected en bloc | 0
lower left pulmonary lobe removed | 0
extubated | 0
spontaneous respiration | 0
SpO2 90% | 0
blood pressure 136/107 mmHg | 0
dyspneic | 5
blood pressure dropped to 65/49 mmHg | 5
dopamine infusion at 5 μg.kg−1.min−1 | 5
rapid fluid infusion | 5
thoracic surgeons notified | 5
blood pressure decreased to 48/37 mmHg | 10
leg elevated | 10
electrocardiogram showed slight inferolateral ST depression | 10
jugular vein engorgement detected | 10
phenylephrine injection | 30
dopamine infusion at 7 μg.kg−1.min−1 | 30
SpO2 decreased to 85% | 30
continuous positive airway pressure of 10 cm H2O | 30
SpO2 increased to 93% | 30
blood pressure dropped to 63/51 mmHg | 105
refractory to high-dose epinephrine and intravascular fluid bolus | 105
dyspnea and tachypnea worsening | 120
intubated | 120
chest X-ray showed haziness in left lung field and enlarged heart with straightened left cardiac border | 120
jugular vein remained distended | 120
Transesophageal Echocardiogram (TEE) performed | 155
moderate pericardial effusion detected | 155
pericardiocentesis attempted | 180
pericardial drainage insufficient | 180
emergency pericardial window operation | 180
600 mL of sanguineous pericardial fluid suctioned | 180
hemodynamics improved dramatically | 180
blood pressure 120/70 mmHg | 180
SpO2 100% | 180
recovered well | 240
outpatient chest X-rays taken during follow-up were clear | 240