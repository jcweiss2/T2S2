76 years old | 0
male | 0
presented to the emergency department | 0
left knee pain | -96
febrile | 0
Glasgow coma scale of 14/15 | 0
heart rate of 125 bpm | 0
polypneic at 25c/min | 0
swelling measuring 15 cm on inner side of left thigh | 0
skin necrosis | 0
inflammatory signs (thigh) | 0
abdomen soft | 0
abdomen not painful | 0
swelling measuring 5 cm in left inguinal region | 0
inflammatory signs (inguinal) | 0
leukocytosis of 30,000E/ml | 0
C-reactive protein of 400 mg/l | 0
computed tomography angiography showing fluid and gas tracking | 0
diagnosis of septic shock | 0
diagnosis of necrotizing fasciitis of left thigh | 0
diagnosis of necrotizing fasciitis of abdominal wall | 0
operation under general anesthesia | 0
hypotension | 0
tachycardia of 150 bpm | 0
high doses of catecholamine | 0
incision in left inner thigh | 0
drainage of 100 milliliters of pus | 0
dissection into quadriceps muscle plains | 0
drainage of 200 milliliters of pus | 0
necrotic debris excised | 0
incision in left inguinal region | 0
dissection into muscle plains | 0
abdominal midline incision | 0
discovery of 5 cm tumor in sigmoid | 0
tumor perforated in retroperitoneum | 0
tumor unresectable | 0
colostomy on left flank | 0
biopsy of tumor | 0
pathological examination showing well-differentiated Lieberkuhnian adenocarcinoma | 0
bacteriological examination showing E. coli multi-drug-sensitive | 0
negative anaerobic culture | 0
septic shock | 0
aggressive debridement of necrotic tissues | 0
high doses of intravenous antibiotics | 0
intensive care support | 0
deceased | 24
