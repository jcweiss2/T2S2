75 years old | 0
    Japanese | 0
    man | 0
    transferred from a local hospital to our intensive care unit | 0
    necrotizing pancreatitis | 0
    smoked 40 cigarettes per day for 50 years | -403200
    old anterior myocardial infarction | 0
    treated with antibiotics | 0
    endoscopic catheter drainage of pancreatic necrosis | 0
    day 8 of admission | 192
    suddenly presented with bradycardia | 192
    suddenly presented with dyspnea | 192
    body temperature of 38.2°C | 192
    blood pressure of 74/52 mmHg | 192
    pulse rate of 50 beats per minute | 192
    oxygen saturation of 91% on 5 L/min oxygen | 192
    elevated white blood cell count (10,900 /μL) | 192
    elevated C-reactive protein level (12.8 mg/dL) | 192
    elevated presepsin level (1,342 pg/mL) | 192
    presence of sepsis | 192
    elevated fibrin degradation products (45.8 μg/mL) | 192
    high prothrombin time-international normalized ratio (1.41) | 192
    low AT activity (49%) | 192
    coagulation disorder | 192
    platelet count within the normal limit | 192
    new-onset ST elevation in inferior leads | 192
    complete atrioventricular block | 192
    reduced left ventricular ejection fraction of 25% | 192
    local hypokinesia in the inferior wall | 192
    local dyskinesia in the anterior wall | 192
    acute inferior myocardial infarction | 192
    old anterior myocardial infarction | 192
    cardiogenic-septic shock | 192
    septic disseminated intravascular coagulation (DIC) | 192
    inserted an intra-aortic balloon pump (IABP) | 192
    inserted a temporary pacemaker | 192
    coronary angiography revealed sub-occlusion of the proximal right coronary artery (RCA) | 192
    started emergent PCI for the RCA | 192
    administered dual antiplatelet agents (200 mg of aspirin and 20 mg of prasugrel) | 192
    administered a bolus of 8,000 units of UFH | 192
    IVUS showed a hypoechoic plaque with deep ultrasound attenuation | 192
    vulnerable plaque at the culprit lesion without visible thrombus | 192
    3.0-mm balloon dilatation | 192
    thrombolysis in myocardial infarction grade 3 flow | 192
    culprit lesion became reoccluded | 192
    preparing stent implantation | 192
    repeat IVUS detected a large build-up of lobulated hypoechoic mobile masses | 192
    fresh thrombi | 192
    aspirated some small red thrombi using a 7-F aspiration catheter | 192
    thrombi remained | 192
    blood flow was not improved | 192
    activated clotting time (ACT) was insufficient at 248 seconds | 192
    used 16,000 units of UFH in total | 192
    suspicion of the presence of HR | 192
    low plasma AT activity | 192
    acquired AT deficiency caused by septic DIC | 192
    administered 2,400 units of AT gamma | 192
    administered additional 5,000 units of UFH | 192
    ACT increased to 364 seconds | 192
    amount of intravascular thrombi decreased | 192
    occluded lesion recanalized | 192
    implanted a drug-eluting stent | 192
    completed PCI without subsequent thrombus formation | 192
    plasma AT activity had increased to 74% | 192
    platelet count did not decrease after PCI | 192
    heparin/platelet factor 4 antibody was not detected | 192
    hemodynamic status was markedly stabilized after the revascularization | 192
    IABP and temporary pacemaker were removed two days after PCI | 216
    required prolonged intensive treatment against refractory pancreatitis | 192
    died due to sepsis on day 45 of admission | 1080
    