74 years old | 0
white | 0
female | 0
admitted to the Emergency Department | 0
low-grade fever | -48
dry cough | -48
shortness of breath | -48
admitted to another hospital for an elective right total knee replacement | -168
pain | -168
redness | -168
swelling | -168
essential hypertension | 0
obesity | 0
myasthenia gravis | 0
osteoarthritis | 0
body temperature of 37.3°C | 0
blood pressure of 121/82 | 0
pulse of 87 beats per minute | 0
respiratory rate of 16 breaths per minute | 0
oxygen saturation of 87% | 0
bilateral rhonchi with rales | 0
patchy air space opacity in the right upper lobe suspicious for pneumonia | 0
rapid nucleic acid amplification test for influenza A and B negative | 0
nasopharyngeal swab specimen obtained | 0
admitted to the airborne-isolation unit | 0
started on broad-spectrum antibiotics with cefepime and levofloxacin | 0
started on 2 L of supplemental oxygen | 0
mild diarrhea | 72
generalized weakness | 72
fatigue | 72
evaluated by Neurology | 72
started on 1 g/kg intravenous immunoglobulin | 72
mild absolute lymphopenia | 0
anemia | 0
pH of 7.46 | 0
pCO2 of 44.6 mmHg | 0
pO2 of 94.7 mmHg | 0
bicarbonate of 31.4 mmol/L | 0
nasopharyngeal swab results came back positive for SARS-CoV-2 | 96
started on oral hydroxychloroquine | 96
started on azithromycin | 96
started on zinc sulfate | 96
started on oral vitamin C | 96
discontinued broad-spectrum antibiotics | 96
SOB worsened rapidly | 144
oxygen requirements went up to 15 L | 144
drowsy | 144
moderate distress | 144
unable to protect the airways | 144
blood pressure of 78/56 mmHg | 144
heart rate of 112 beats per minute | 144
temperature of 38°C | 144
respiratory rate of 28 breaths per minute | 144
bilateral alveolar infiltrates due to pneumonia and interstitial edema consistent with ARDS | 144
intubated | 144
started on pressure-regulated volume-controlled mechanical ventilation | 144
started on norepinephrine | 144
started on colchicine | 144
started on high-dose vitamin C | 168
norepinephrine support stopped | 192
CXR showed significant improvement of the pneumonia and interstitial edema | 240
spontaneous breathing trial with CPAP/PS | 240
tolerated by the patient | 240
pH of 7.49 mmHg | 240
pCO2 of 40.2 mmHg | 240
pO2 of 77.1 mmHg | 240
bicarbonate of 30.2 mmol/L | 240
extubated to 4 L of oxygen with a nasal cannula | 240
breathing status continued to improve | 384
oxygen saturation of 92% | 384
CXR revealed almost complete resolution of the infiltrates | 384
discharged from the hospital | 384