73 years old | 0
female | 0
established renal failure | 0
poor vessels for primary or secondary vascular access | 0
admitted electively | 0
creation of a first-stage brachiobasilic arteriovenous fistula | 0
transferred to haemodialysis | -672
peritonitis | -672
laparotomy | -672
tunnelled jugular central venous catheter | -504
metallic mitral valve replacement | -10080
therapeutic anticoagulation | -10080
hypertension | -10080
haematuria | -10080
diarrhoea | -72
rigours | -72
pain around her line | -72
treatment for presumed catheter-associated bacteraemia | -72
septic | -72
swinging fevers | -72
splinter haemorrhage | -72
new murmur | -72
possible vegetation on her mitral valve | -72
blood cultures positive for Staphylococcus aureus | -72
treatment for endocarditis | -72
antibiotics | -72
responded well to treatment | -24
represented feeling unwell | 672
non-specific symptoms | 672
routine observations normal | 672
blood investigations normal | 672
lactic acidosis | 672
mild lower abdominal pain | 672
fast, uncontrolled atrial fibrillation | 672
arterial blood gas | 672
pH 7.13 | 672
pO2 103 mmHg | 672
pCO2 17.3 mmHg | 672
lactate 13.3 mmol/L | 672
contrast-enhanced CT angiogram | 672
patent celiac and superior mesenteric artery axis | 672
patent portal vein | 672
chronic pyelonephritis | 672
possible inflammation in the gallbladder fossa | 672
inflammatory oedema in Morrison’s pouch | 672
transferred to intensive care unit | 672
resuscitated | 672
intubated | 672
ventilated | 672
haemodynamically stable | 672
metabolic acidosis worsened | 672
arterial lactic acid increased | 672
emergency laparotomy | 696
sero-purulent fluid in Morrison’s pouch | 696
macro-nodular liver | 696
normal gallbladder | 696
stomach, duodenum and pancreas normal | 696
small bowel and colon normal | 696
extensive inflammatory change around the right kidney | 696
nephrectomy | 696
haemofiltered | 700
speedy recovery | 704
arterial lactic acid returned to normal | 704
discharged to the ward | 752
pathology revealed chronic pyelonephritis | 752
sclerosis of the glomeruli | 752
atrophy of the tubules | 752
polymorphs | 752
chronic inflammation | 752
fibrosis of the parenchyma | 752
no evidence of renal stones | 752
hypertensive change in arterioles | 752
final diagnosis of chronic pyelonephritis with peri-renal sepsis | 752
liver biopsy | 752
congestive hepatomegaly | 752