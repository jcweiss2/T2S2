stabs herself in the abdomen with a kitchen knife | -1
admitted to emergency department | 0
blood pressure could not be measured | 0
pulseless electrical activity | 0
body temperature was 35.0 °C | 0
oxygen saturation was 99 % | 0
Glasgow Coma Scale score of 3 | 0
agonal respiration | 0
wound measuring 5 cm on upper abdomen | 0
intra-abdominal fluid collection | 0
emergency thoracotomy | 0.5
aortic cross-clamping | 0.5
open cardiac massage | 0.5
administration of epinephrine | 0.5
temporary return of spontaneous circulation | 1
hemodynamically unstable | 1
laparotomy | 1
injuries to common hepatic and splenic arteries | 1
injuries to pancreas, spleen, and liver | 1
ligation of injured arteries | 1
distal pancreatectomy | 1.5
splenectomy | 1.5
liver sutured | 1.5
administration of norepinephrine | 1.5
second-look surgery | 24
no active bleeding or ischemic change | 24
no vasopressor requirement | 72
abdominal wall closure | 72
enhanced computed tomography scan | 96
disruption of celiac artery | 96
gastroduodenal artery arising from superior mesenteric artery | 96
gastroscopy | 216
patchy mucosal necrosis on gastric upper body | 216
conservative treatment | 216
fever of 39 °C | 552
pain in stomach | 552
white blood cell count of 34,000/mm3 | 552
C reactive protein of 13.4 mg/dL | 552
CT scan | 552
air in gastric wall | 552
intra-abdominal free air | 552
gastric necrosis | 552
emergency surgery | 552
total gastrectomy with Roux-en-Y reconstruction | 552
histological findings of stomach | 552
diffuse necrotic changes | 552
inflammatory cell infiltrations | 552
no evidence of invasive fungal infection | 552
leakage on duodenal stump | 696
continuous tube drainage | 696
sepsis due to multidrug-resistant Pseudomonas aeruginosa infection | 1680
disseminated intravascular coagulation | 1680
death | 1680