44 years old | 0
male | 0
admitted to the hospital | 0
pleuritic chest pain | 0
fever | 0
chills | 0
night sweats | 0
persistent chest pain | 0
tachycardia | 0
oxygen saturation of 92% | 0
mild distress | 0
distant heart sounds | 0
no pericardial rubs | 0
oral temperature of 97.9°F | 0
blood pressure of 110/71 mm Hg | 0
pulsus paradoxus not present | 0
pulmonary sarcoidosis | -336
EBUS bronchoscopy | -336
mediastinal and hilar lymphadenopathy | -336
chest computed tomography | -336
noncaseating granulomas | -336
essential hypertension | -10080
smoking denied | 0
alcohol use denied | 0
illicit drug use denied | 0
prior international travel denied | 0
pet ownership denied | 0
chest x-ray | -5184
scattered pulmonary nodules | -5184
comprehensive chest CT | -5184
small scattered pulmonary nodules | -5184
COVID-19 pneumonia | 0
acute pericarditis | 0
pulmonary embolism | 0
myocarditis | 0
acute coronary syndrome | 0
electrocardiogram | 0
diffuse ST-segment elevations | 0
PR depression | 0
serial negative troponin | 0
D-dimer >250 ng/mL | 0
C-reactive protein of 204.5 mg/L | 0
sedimentation rate of 65 mm/h | 0
chest CT with pulmonary angiography | 0
no pulmonary embolism | 0
circumferential pericardial effusion | 0
worsening of multiple diffuse pulmonary nodules | 0
negative blood cultures | 0
transthoracic echocardiogram | 0
preserved left ventricular ejection fraction | 0
moderate-size circumferential pericardial effusion | 0
early diastolic right ventricular collapse | 0
significant variation in mitral inflow E velocity | 0
plethoric inferior vena cava | 0
supplemental oxygen | 0
oral analgesia | 0
echocardiography-guided pericardiocentesis | 2
drainage of 250 mL of purulent material | 2
admitted to the intensive care unit | 2
broad spectrum antibiotics | 2
intravenous piperacillin/tazobactam | 2
intravenous vancomycin | 2
pericardial drain | 2
pericardial drain removal | 128
worsening of left pleural effusion | 96
left thoracocentesis | 96
left chest tube placement | 96
intrapleural thrombolysis | 96
exudative process | 96
fluid cultures grew Actinomyces odontolyticus | 96
antibiotics de-escalated | 96
intravenous ampicillin-sulbactam | 96
chest tube removal | 168
pericardial effusion recurred | 240
no clinical or echocardiographic tamponade | 240
pericardial window via left anterior thoracotomy | 312
inflammatory markers improved | 360
discharged | 360
CRP of 19 mg/L | 360
sedimentation rate of 40 mm/h | 360
no recurrence of acute pericarditis | 360