74 years old | 0
female | 0
ulcerative colitis | -6720
colectomy | -6720
ileostomy | -6720
hypertension | -6720
admitted to the hospital | 0
fatigue | 0
myalgia | 0
confusion | 0
temperature of 100°F | 0
blood pressure of 108/60 mmHg | 0
heart rate of 106 bpm | 0
respiratory rate of 20 breaths per minute | 0
disoriented to the surrounding environment | 0
normal S1 and S2 without murmurs, gallops or rubs | 0
decreased breath sounds on lung bases without crackles or rales | 0
sodium of 128 | 0
creatinine of 1.21 | 0
elevated lactate at 3.0 | 0
urinalysis suggestive of urinary tract infection (UTI) | 0
white blood cell count of 8.8 | 0
hemoglobin of 15.1 | 0
platelet count of 131 | 0
CT of the brain unremarkable | 0
chest X-ray unremarkable | 0
resuscitated with intravenous fluid | 0
started on IV ceftriaxone | 0
admitted for treatment of sepsis | 0
discharged | 72
returned to the ED | 96
complaint of significant weakness | 96
inability to ambulate | 96
elevated temperature of 103°F | 96
heart rate of 115 bpm | 96
blood pressure of 90/65 mmHg | 96
respiratory rate of 24 breaths per minute | 96
normal mental status | 96
white blood cell count of 3.31 | 96
hemoglobin of 13.2 | 96
platelet count of 60 | 96
lactic acid of 5.4 | 96
AST of 237 | 96
ALT of 189 | 96
alkaline phosphatase of 146 | 96
Chest X-ray showed right middle lobe infiltrates | 96
started on vancomycin and piperacillin-tazobactam | 96
admitted to the medical floor | 96
worsening respiratory status | 120
noninvasive mechanical ventilation | 120
transferred to the medical intensive care unit | 120
bilateral pleural effusions on CT of the chest | 120
thoracentesis | 120
removal of 750cc of exudative fluid | 120
progressively hypoxemic | 120
serial chest X-rays showing bilateral interstitial infiltrates | 120
intubation | 120
fever persisted | 120
decline in her state | 120
multiple blood, sputum, urine, and stool cultures negative | 120
white blood cell count of 1.4 | 144
hemoglobin of 8.5 | 144
platelet count of 45 | 144
worsening kidney functions tests | 144
creatinine of 2.1 | 144
BUN of 65 | 144
liver transaminases continued to rise | 144
jaundice worsened | 144
coagulopathy | 144
elevated international normalized ratio (INR) at 8 | 144
acute liver injury (ALI) | 144
Factor V and factor VIII activity assays normal | 144
ruled out disseminated intravascular coagulopathy (DIC) | 144
abdominal ultrasound unremarkable | 144
MRI of the liver and pancreas unremarkable | 144
elevated LDH at 1367 | 144
elevated triglycerides at 808 | 144
fibrinogen of 240 | 144
elevated ferritin at 40,000 | 144
suspected HLH | 144
bone marrow biopsy | 144
normocellular marrow with myeloid predominance | 144
mild granulocyte atypia | 144
increased histiocytes | 144
CD163 immunostaining of the core biopsy | 144
markedly increased histiocytes with some cells showing ingested cellular material | 144
started on an 8-week-regimen of dexamethasone and etoposide | 144
improvement of her clinical status | 168
cell counts improved | 168
liver functions improved | 168
viral serologies obtained | 168
negative for human immunodeficiency virus (HIV) | 168
negative for cytomegalovirus (CMV) | 168
negative for Herpes simplex virus (HSV) type 1 and 2 | 168
negative for Epstein-Barr virus (EBV) | 168
negative for hepatitis B virus | 168
negative for hepatitis C virus | 168
antinuclear antibody negative | 168
double-stranded DNA antibody negative | 168
rheumatoid factor negative | 168
autoimmune hepatitis workup negative | 168
hereditary hemochromatosis ruled out | 168
DNA assay for C282Y, H63D, and S65C loci of the gene HFE showed no mutations | 168
diagnosed with HLH | 168
met 5 out of the 8 criteria | 168
fever | 168
cytopenia of 2 cell lines | 168
elevated ferritin>500 ng/mL | 168
elevated fasting triglyceride >265 mg/dL | 168
hemophagocytosis in bone marrow | 168
respiratory status improved | 216
weaned off mechanical ventilation | 216
blood counts improved dramatically | 216
normalization of liver enzymes | 216
readmitted to the hospital | 744
persistent confusion | 744
diagnosed with HLH with central nervous system involvement | 744
started on intrathecal methotrexate | 744
no improvement in her symptoms | 744
goals of care changed to comfort care | 744
passed away | 768