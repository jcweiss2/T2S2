66 years old | 0
male | 0
history of Billroth II gastrectomy for peptic ulcer disease | -302400
history of open cholecystectomy | -87600
presented to the emergency department | 0
diffuse abdominal pain | 0
vomiting | 0
diarrhea | 0
admitted receiving nonsteroidal anti-inflammatory drugs | 0
admitted receiving colchicine | 0
persisting gout crisis | 0
diffuse articular pain | 0
afebrile | 0
mild tenderness to deep palpation in all four abdominal quadrants | 0
rectal examination revealed enlarged prostate | 0
marked leukocytosis (48,000/mm3) | 0
INR of 2.5 | 0
C-reactive protein of 48 mg/l | 0
arterial blood gas pH 7.21 | 0
base excess of 13.6 mEq/l | 0
pCO2 of 33 mmHg | 0
judged as not having acute abdominal disease | 0
plain abdominal X-ray showed no pathology | 0
ultrasound showed simple left renal cyst | 0
computed tomography scan showed dilatation and edema of jejunal loops | 0
computed tomography scan showed minimal free fluid in peritoneal space | 0
radiology report suggested localized peritonitis | 0
developed respiratory failure | 2
required intubation | 2
required mechanical ventilation | 2
became severely hypotensive (60/40 mmHg) | 2
became oliguric | 2
initiated inotropic support | 2
noted macroscopic hematuria | 2
possibility of intra-abdominal collection not ruled out | 2
no other source of septic shock identified | 2
emergency explorative laparotomy decided | 2
laparotomy found no anastomotic leak | 2
laparotomy found no source of abdominal sepsis | 2
continued multiorgan failure | 16
died | 16
colchicine overdose diagnosed postmortem | 16
