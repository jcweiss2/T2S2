69 years old | 0
woman | 0
presented to the emergency department | 0
high-grade fever | -72
pleuritic right lower chest pain | -72
cough | -72
elevated temperature of 38.8°C | 0
bibasilar crackles | 0
lower extremity edema | 0
grade 3 holosystolic apical murmur | 0
mitral valve regurgitation | 0
long-term venous access port | -26208
recurrent transfusion-dependent anemia | -26208
hemoglobin 12.1 g/dL | 0
white blood cell count 15.1×103/µL | 0
absolute neutrophil count 13.2×103/µL | 0
b-type natriuretic peptide 788 pg/mL | 0
chest radiography changes consistent with congestive heart failure | 0
electrocardiography showed left bundle branch pattern | 0
blood cultures positive for Corynebacterium CDC group G | 0
gram stain positive for gram positive rods | 0
transthoracic echocardiography demonstrated moderate mitral valve regurgitation | 0
thickened anterior mitral leaflet suggesting vegetations | 0
pulmonary artery systolic pressure of 84 mmHg | 0
echocardiogram one year prior without mitral valve thickening | -8760
diagnosed with bacterial IE secondary to Corynebacterium CDC group G | 0
involvement of the mitral valve | 0
penicillin allergy | 0
treated with intravenous vancomycin | 0
treated with clindamycin | 0
6-week course of antibiotics | 0
chronic implanted venous access port removed | 0
discharged to extended care facility | 0
readmitted due to sudden onset shortness of breath | 72
hypoxic | 72
white blood cell count elevated to 18×103/µL | 72
vancomycin therapy continued | 72
repeat transthoracic echocardiography showed severe mitral valve regurgitation | 72
large and mobile vegetation on the mitral valve | 72
mitral valve replacement with 27-mm Edwards-Carpentier pericardial valve | 72
coronary artery bypass grafting surgery | 72
reverse saphenous vein graft to the distal right coronary artery | 72
native mitral valve leaflet pathology revealed endocarditis | 72
fibrinopurulent exudate | 72
granulation tissue | 72
cultures positive for diphtheroids | 72
post-operative oliguric acute renal failure | 72
respiratory failure requiring mechanical ventilation | 72
urinary tract infection with vancomycin resistant enterococcus | 72
vancomycin discontinued | 72
daptomycin therapy started | 72
worsening congestive heart failure | 168
transesophageal echocardiogram on day 17 of re-admission | 408
severe mitral valve regurgitation | 408
well-seeded mitral valve annular plane | 408
echo densities on the mitral valve leaflets | 408
recurrent endocarditis of prosthetic valve | 408
antibiotic therapy broadened with doxycycline | 408
antibiotic therapy broadened with aztreonam | 408
antibiotic therapy broadened with anidulafungin | 408
daptomycin continued | 408
porcine valve replaced with mechanical St. Jude’s prosthesis | 408
intraoperative transesophageal echocardiogram confirmed well-functioning prosthetic mitral valve | 408
bioprosthetic mitral valve pathology showed fibrous and fibro-inflammatory tissue | 408
cultures remained negative | 408
limb ischemia | 504
bleeding through orifices and lines | 504
elevation of partial thromboplastin time | 504
elevation of prothrombin time | 504
disseminated intravascular coagulation | 504
multi-organ failure | 504
expired | 504
prior blood cultures positive for diphtheroids 4 months prior | -2880
line-associated bacteremia not entertained | -2880
identification not done | -2880
