43 years old | 0
male | 0
admitted to the hospital | 0
upper abdominal pain | -24
colic | -24
vomiting | -24
diarrhea | -24
history of similar attacks | -24
afebrile | 0
hemodynamically stable | 0
tender right upper abdominal part | 0
positive Murphy's sign | 0
leucocytosis | 0
liver function tests normal | 0
electrolytes normal | 0
gall bladder stone | 0
acute cholecystitis | 0
treated with intravenous fluids | 0
treated with ceftriaxone | 0
treated with metronidazole | 0
treated with dalteparin | 0
laparoscopic cholecystectomy | 6
edematous gall bladder | 6
single stone | 6
adhesions | 6
intra-abdominal pressure 12-15 mmHg | 6
histopathology report showed acute cholecystitis | 6
histopathology report showed chronic cholecystitis | 6
recovered well | 48
scheduled to be discharged | 48
new severe epigastric pain | 48
severe leucocytosis | 48
partial obstruction at the origin of the SMA | 48
ischemia of the small bowel | 48
obstruction and dilatation of the proximal part of the small bowel | 48
abdominal exploration | 72
ischemic terminal ileum | 72
good pulsation of the SMA | 72
resection and anastomosis of the ileum | 72
Bogota bag closure of the abdomen | 72
transferred to the SICU | 72
fully heparinized | 72
intubated | 72
sedated | 72
ventilated | 72
second look laparotomy | 96
viable healthy bowel | 96
no leakage at the anastomosis site | 96
abdominal wall closed | 96
heparinization resumed | 102
started on total parental nutrition | 102
normal echocardiogram | 102
no deep venous thrombus | 102
sinus rhythm | 102
abdominal distension increased | 288
elevation of the IAP to 24 mmHg | 288
hemoglobin dropped to 6.3 g/dl | 288
received blood and blood products | 288
abdominal collections | 312
condition deteriorated | 336
abdomen more distended | 336
required full ventilatory support | 336
oliguric | 336
elevation of the IAP to 25 mmHg | 336
diagnosed as ACS | 336
decompressive laparotomy | 336
old and partially hemolysed blood-stained fluid collection drained | 336
abdomen closed by using a bagota bag | 336
unstable and needed inotropic support | 336
highly febrile | 360
septic shock | 360
renal failure | 360
started on renal replacement therapy | 360
asystole | 384
died | 384