55 years old | 0
female | 0
admitted to the hospital | 0
abdominal distress | 0
2 kidney transplantations | -10080
IgA nephropathy | -10080
first allograft lost due to chronic allograft rejection | -10080
current allograft functioning with estimated glomerular filtration rate of approximately 60 ml/min per 1.73 m2 | 0
computed tomographic scan revealed free intra-abdominal air | 0
sigma perforation | 0
sigma resection | 0
protective ileostomy | 0
burst abdomen | 24
surgical intervention for burst abdomen | 24
presumed peritonitis | 48
surgical intervention for presumed peritonitis | 48
fever | 72
respiratory insufficiency | 72
hemodynamic compromise | 72
mechanical ventilation | 72
norepinephrine | 72
antibiotic therapy intensified | 72
vitamin C administration | 72
vitamin B1 administration | 72
urine output decline | 96
plasma creatinine increase | 96
tubular proteinuria | 96
urine microscopy | 96
sonography excluded obstructive uropathy | 96
vascular resistance indices of the kidney allograft within normal range | 96
continuous renal replacement therapy initiated | 120
kidney allograft biopsy | 120
acute tubular injury | 120
oxalate nephropathy | 120
vitamin C discontinued | 120
citrate-based renal replacement therapy | 120
urinary output restored | 168
continuous renal replacement therapy terminated | 168
second episode of acute kidney injury | 720
kidney allograft function recovered | 8760
estimated glomerular filtration rate of approximately 45-50 ml/min per 1.73 m2 | 8760
discharged | 720