61 years old | 0
male | 0
dyspnea | -120
fever | -120
diagnosed with COVID-19 | -120
hospitalized | -120
thoracic computed tomography | -120
multiple infiltrates in both lungs | -120
treatment with hydroxychloroquine | -120
treatment with azithromycin | -120
treatment with favipiravir | -120
admitted to ICU | -114
tachypnea | -114
high level of oxygen demand | -114
moderate respiratory distress | -114
oxyhemoglobin saturation of 91% | -114
treated with tocilizumab | -114
CRS | -114
severe lymphopenia | -114
hyperferritinemia | -114
prone position | -114
high-flow oxygen support | -114
rapidly progressed to acute hypoxemic respiratory failure | -112
second dose of tocilizumab | -112
intubated | -112
worsening hypoxemia | -112
accessory muscle use | -112
paradoxical abdominal respiration | -112
central venous catheter | -112
mechanical ventilation support | -112
extubated | -96
complained of right shoulder and chest pain | -24
pain radiating to the right arm | -24
exacerbated by sneezing | -24
exacerbated by coughing | -24
exacerbated by deep breathing | -24
exacerbated by movements of the right shoulder and torso | -24
afebrile | -24
bilateral upper extremity muscle strength normal | -24
glenohumeral joint range of motion normal | -24
active and passive movements of the right shoulder extremely painful | -24
redness around the right parasternal region | -24
warmth around the right parasternal region | -24
swelling around the right parasternal region | -24
pain in a referred distribution | -24
mildly elevated serum C-reactive protein | -24
normal leukocyte count | -24
moderate lymphopenia | -24
diagnosed with Tietze syndrome | -24
treated with paracetamol | -24
pain progressively increased | -18
pain spread into the neck | -18
treated with diclofenac | -18
treated with tramadol | -18
oxygen-dependent | -18
treated with methylprednisolone | -18
shoulder and chest pain increased | -18
sternoclavicular joint swollen | -18
sternoclavicular joint red | -18
sternoclavicular joint tender | -18
fluid collection in the right sternoclavicular joint | -18
extension into the chest cavity | -18
chest wall abscess | -18
inflammatory changes | -18
central avascular area within the abscess | -18
CT-guided fine needle aspiration | -18
purulent liquid | -18
Gram stain showed numerous polymorphonuclear leucocytes | -18
acid-fast stain negative | -18
culture of the liquid revealed methicillin-sensitive Staphylococcus aureus | -18
beta-lactam allergy | -18
treated with linezolid | -18
responded well to therapy | -12
discharged home | -12
treated with clindamycin | -12
CT and MRI performed at one month of follow-up | 720
decrease in the diameter and content of the abscess | 720