54 years old | 0
male | 0
admitted to the hospital | 0
pre-syncope | 0
syncope | 0
left-sided chest tightness | 0
generalized fatigue | -672
weight loss | -672
diffuse erythematous rash | 0
blood pressure of 96/60 mm Hg | 0
unremarkable cardiac examination | 0
unremarkable respiratory examination | 0
normal sinus rhythm | 0
raised troponin concentration | 0
eosinophil count of 7.6 × 10^9/l | 0
referred to cardiology | 0
myocarditis | 0
cardiac magnetic resonance imaging | 24
eosinophilic myocarditis | 24
coronary angiography | 24
no evidence of coronary artery disease | 24
skin biopsy | 48
cardiac biopsy | 48
edoxaban | 72
prednisolone | 72
discharged | 72
missed appointment | 1344
presented to cardiology clinic | 1344
neck swelling | 1344
urgently admitted to hospital | 1344
rise in eosinophil count | 1344
increase dose of prednisolone | 1344
computed tomography of neck | 1344
lymphadenopathy | 1344
T-cell lymphoma | 1344
cyclophosphamide | 1344
sepsis | 1400
cholecystitis | 1400
new onset of seizures | 1400
reduction in consciousness | 1400
Glasgow Coma Scale of 9/15 | 1400
head CT | 1400
multiple bilateral acute infarctions | 1400
transferred to intensive care unit | 1400
history of hepatitis B | 0
history of asthma | 0
history of intravenous drug use | 0
history of excessive use of alcohol | 0
ischemic stroke | 1400
reduced GCS score | 1400
seizures | 1400
intracranial bleeding | 1400
malignancy | 1400
intracerebral infection | 1400
diffuse subendocardial late gadolinium enhancement | 1400
mild LV systolic impairment | 1400
eczematous changes | 1400
bone marrow biopsy | 1400
axillary lymph node biopsy | 1400
infarcts involving frontal, parietal, and left temporo-occipital regions | 1400
apical tear | 1400
intramural myocardial tear | 1400
small apical cavity | 1400
diastolic flow in apical cavity | 1400
systolic flow out of apical cavity | 1400
cyclophosphamide therapy | 1400
partial response | 1400
reduction of eosinophil count | 1400
palliation | 1440