32 years old | 0
primigravida | 0
dichorionic twin pregnancy | 0
admitted to emergency department | 0
preterm rupture of membranes of the first fetus | 0
spontaneous dichorionic twin pregnancy | 0
blood type O Rh-positive | 0
ultrasound revealed two viable twins | 0
normal growth for gestational age | 0
oligohydramnios of the first fetus | 0
normal cervical length | 0
subserous uterine fibroid | 0
spontaneous onset of labor | -168
female baby weighing 340 g | -168
vaginal delivery | -168
fetal death occurred within 1 h | -168
histopathological examination showed multi-organic congestion | -168
uterine contractions ceased | -168
cervix reconstituted | -168
no signs of chorioamnionitis | -168
amniotic membrane of the second twin intact | -168
ultrasonography showed healthy remaining fetus | -168
umbilical cord of the first fetus ligated | 0
placenta left inside the uterus | 0
cervical cultures taken | 0
perineum and vagina disinfected with chlorhexidine | 0
patient remained in hospital | 0
treated with bed rest | 0
low-molecular-weight heparin | 0
broad-spectrum antibiotics | 0
ampicillin | 0
gentamycin | 0
amoxicillin | 0
continuous monitoring | 0
clinical assessment | 0
laboratory tests | 0
no signs of infection | 0
serial ultrasonography revealed normal fetal growth | 0
wellbeing of the second twin | 0
digital vaginal examinations avoided | 0
antenatal corticosteroids administered | -96
betamethasone | -96
urgent cesarean section due to breech presentation | 24
spontaneous labor | 24
female neonate weighing 685 g | 24
Apgar scores 1/8/9 | 24
full resuscitation | 24
immediate life-support intervention | 24
admitted to Neonatal Intensive Care Unit | 24
extreme prematurity | 24
extreme low birth weight | 24
Hyaline membrane disease | 24
patent ductus arteriosus | 24
satisfactory evolution | 24
spontaneous respiration at one month | 24
discharged 90 days after birth | 24
postpartum sepsis due to endometritis | 24
admitted to Intensive Care Unit | 24
discharged 12 days after surgery | 24
no complications | 24
normal cognitive development at 15th month | 24
normal neurological development at 15th month | 24
low weight | 24
deficient physical development for age | 24
patent ductus arteriosus maintained | 24
