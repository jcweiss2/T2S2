61 years old | 0
female | 0
non-smoking | 0
veteran | 0
hypertension | -672
chronic cough | -168
dyspnea | -168
weight loss | -168
nausea | -72
vomiting | -72
cachexia | 0
scleral icterus | 0
jaundice | 0
dry mucous membranes | 0
decreased breath sounds | 0
tachycardia | 0
hypotension | 0
hyponatremia | 0
elevated alkaline phosphatase | 0
elevated total bilirubin | 0
elevated aspartate aminotransferase | 0
elevated alanine aminotransferase | 0
pulmonary parenchymal nodules | 0
pleural effusion | 0
pancreatic head mass | 0
biliary ductal dilation | 0
lung adenocarcinoma | 0
brain metastases | 0
radiation therapy | 24
chemotherapy | 24
biliary stenting | 24
biopsy of lung mass | 24
biopsy of pancreatic head | 24
high nuclear pleomorphism | 24
prominent nuclei | 24
positive TTF-1 staining | 24
positive CK-7 staining | 24
negative p63 staining | 24
severe pneumonia | 168
sepsis | 168
death | 168