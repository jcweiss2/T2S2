64 years old | 0
female | 0
elective radical total gastrectomy | 0
feeding jejunostomy | 0
poorly differentiated T1 gastric carcinoma | 0
hypertension | -672
anaemia | -672
antihypertensive medication | -672
jejunostomy feeds commenced | 24
routine post-operative contrast CT scan | 48
bilateral pleural effusions | 48
multiple vomits | 96
not opened bowels since procedure | 96
tachycardic | 96
febrile | 96
dyspnoeic | 96
mildly tender abdomen | 96
cool peripheries | 96
pH 7.45 | 96
Lactate 4.2 mmol/L | 96
white cell count 1.9 × 10^9/L | 96
C-reactive protein 456 mg/L | 96
septic workup | 96
repeat CT chest abdomen pelvis | 96
broad spectrum antibiotics | 96
suspected aspiration pneumonia | 96
dilated roux loop | 96
obstruction | 96
distended caecum | 96
ascending colon | 96
caecal volvulus | 96
urgent exploratory laparotomy | 120
grossly distended caecal volvulus | 120
compressing feeding jejunostomy | 120
obstructing small bowel | 120
right hemicolectomy | 120
jejunostomy un-kinked | 120
small bowel viability confirmed | 120
feeding tube removed | 120
small bowel defect repaired | 120
bacteraemia | 144
intravenous antibiotics | 144
tracheostomy | 168
ARDS | 168
pericardial effusion | 168
pleural effusions | 168
full recovery | 720
ischaemic changes | 720 
histology of resected colon | 720