21 years old | 0
primigravida | 0
16 weeks gestation | 0
asthma | 0
depression | 0
anxiety | 0
presented to urgent care clinic | -240
suspected streptococcal pharyngitis | -240
discharged on oral Amoxicillin | -240
completed Amoxicillin | -240
presented to ED | -168
fever | -168
sore throat | -168
discharged home | -168
broke out in a rash | -168
presented to OSH ED | -168
fever 104°F | -168
body aches | -168
dry cough | -168
rash | -168
prenatal vitamin supplement | 0
temperature 103.8°F | 0
blood pressure 109/57 mmHg | 0
pulse 114 beats per minute | 0
respiratory rate 18 breaths per minute | 0
oxygen saturation 98% | 0
erythematous plaques | 0
indurated plaques | 0
subtle scaling | 0
vesicles on hands | 0
vesicles on feet | 0
vesicles on mouth | 0
ulcers in hard palate | 0
lactate 2.6 | 0
white blood cell count 3.3 k/ul | 0
hemoglobin 8.3 g/dl | 0
platelets 157 k/ul | 0
spherocytes on blood smear | 0
chest x-ray unremarkable | 0
intravenous fluids | 0
IV antibiotics | 0
suspected sepsis | 0
negative blood cultures | 24
negative throat culture | 24
negative MRSA culture | 24
met SIRS criteria | 24
tachycardic | 24
tachypneic | 24
transferred to our facility | 24
febrile | 72
tachycardic | 72
borderline hypotensive | 72
started on high-flow nasal cannula | 72
IV azithromycin | 72
IV cefepime | 72
IV vancomycin | 72
oral acyclovir | 72
switched to IV acyclovir | 72
persistent fevers | 72
tachycardia | 72
tachypnea | 72
acutely dyspneic | 96
hypoxic 88% | 96
CXR bilateral pleural effusions | 96
multifocal pneumonia | 96
pulmonary edema | 96
CT chest bilateral airspace disease | 96
continued antibiotics | 96
negative infectious workup | 96
endotracheal intubation | 96
mechanical ventilation | 96
hemoglobin decreased | 96
leukopenia 2.6 K/dL | 96
thrombocytopenia 119 K/dL | 96
lymphopenia | 96
negative hemolysis | 96
positive Coombs test | 96
elevated LDH | 96
normal haptoglobin | 96
positive ANA 1:640 | 96
anti-RNP 113 | 96
anti-Smith 103 | 96
complement C3 26 | 96
complement C4 <8 | 96
negative autoantibodies | 96
interface dermatitis | 96
vacuo-lar changes | 96
vascular damage | 96
BAL alveolar hemorrhage | 96
Candida albicans in BAL | 96
negative viral panels | 96
negative bacterial panels | 96
proteinuria 1.83 g/24h | 96
no lupus nephritis | 96
IV methylprednisolone | 96
plasmapheresis | 96
multi-specialty collaboration | 96
cyclophosphamide consented | 96
high fever | 120
hypotension | 120
tachycardia | 120
candidemia | 120
treated with fluconazole | 120
bilateral cotton wool spots | 120
extubated | 120
cyclophosphamide 500 mg | 120
acute abdominal pain | 192
lipase 1688 | 192
amylase 560 | 192
alkaline phosphatase 55 IU/L | 192
total protein 5.2 g/dL | 192
total bilirubin 1.0 md/dL | 192
albumin 2.6 g/dL | 192
CT confirmed acute pancreatitis | 192
discharged on hydroxychloroquine | 216
prednisone taper | 216
preterm premature rupture of membranes | 672
spontaneous labor | 672
magnesium sulfate | 672
delivered healthy baby | 672
