65 years old | 0
woman | 0
admitted to the hospital | 0
worsening respiratory distress | 0
low back pain | 0
transferred to the intensive care unit | 24
took bisphosphonate | -24
osteoporosis | -24
blood pressure 132/85 mmHg | 0
pulse rate 145/min | 0
hematocrit 39% | 0
white-cell count 10,300/mm3 | 0
serum urea nitrogen 58 mg/dl | 0
creatinine 1.85 mg/dl | 0
serum sodium 128 mEq/L | 0
potassium 5 mEq/L | 0
chloride 101 mEq/L | 0
lactate dehydrogenase 345 | 0
serum glutamic oxaloacetic transaminase 90 U/L | 0
creatine kinase 422 U/L | 0
bilirubin 3.07 mg/dl |3 0
abnormal coagulation profile | 0
disseminated intravascular coagulation | 0
contrast-enhanced computed tomography of the abdomen | 0
hypodense zone of the renal cortex | 0
hyperdense medulla | 0
no excretion of contrast media into the collecting system | 0
hemodialysis | 24
anticoagulation | 24
supportive measures | 24
condition deteriorated | 168
died | 168
