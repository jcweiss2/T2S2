18 years old | 0
male | 0
admitted to the hospital | 0
fever | 0
scrotal pain | 0
tachycardia | 0
hypotension | 0
broad-spectrum antibiotics | 0
vancomycin | 0
Zosyn | 0
switched to meropenem | 0
acute kidney injury | 0
fever persisted | 0
no source of infection found | 0
stopping all antibiotics | 0
macular rash | -120
rash progressed | -96
axillary area involved | -96
chest involved | -96
head involved | -96
neck involved | -96
abdomen involved | -96
decline of mental status | -96
worsening of skin lesions | -96
bullae and vesicles | -96
rash became pustular | -72
high grade fever | -72
pulse steroids | -72
fever subsided | -69
rash improved | -69
sloughing decreased | -69
acute kidney injury resolved | -69
taper in steroids | -69
skin biopsy | -69
intra- and subcorneal spongiform | -69
superficial, interstitial, mid-dermal infiltrate rich in neutrophils | -69
dermal edema | -69
DRESS | -69
GPP | -69
PAN typical rash | -69
Steven Johnson syndrome | -69
leukocytoclastic vasculitis | -69
subcorneal pustular dermatosis | -69
cutaneous candidiasis | -69
fever and leukocytosis | -672
acute kidney injury | -672
Zosyn | -672
meropenem | -672
re-challenged with meropenem and vancomycin | -672
no reaction | -672
PAN | -672
multiple prior admissions | -672
septic shock | -1344