41 years old | 0
female | 0
admitted to the hospital | 0
acute stabbing upper abdominal pain | -48
radiating to the scapula | -48
no vomiting | -48
no reflux | -48
no dysphagia | -48
normal bowel habits | -48
weight 70 kg | 0
body mass index (BMI) 26.35 kg/m2 | 0
gained 2 kg during pregnancy | 0
BMI before conception 25.6 kg/m2 | -9360
laparoscopic gastric band insertion | -9360
third pregnancy | 0
one missed abortion | -9360
one previous caesarean delivery | -9360
obstetrical scans at 13th week | -728
no pathologies detected | -728
obstetrical scans at 19th week | -560
no pathologies detected | -560
hyperemesis gravidarum | -728
mild constipation | -728
abdominal pain at 18th week | -504
lower abdomen pain | -504
left lumbal region pain | -504
umbilical region pain | -504
appendicitis suspected | -504
admitted to surgery department | -504
C-reactive protein (CRP) 23 mg/l | -504
C-reactive protein (CRP) 40 mg/l | -502
diagnosis of appendicitis excluded | -502
discharged from hospital | -502
referred to perinatology center | -502
no further medical attention | -502
blood pressure 90/62 mmHg | 0
pulse rate 112 bpm | 0
positive Blumberg sign | 0
leukocytosis 22.89 x 10^9/l | 0
CRP 289.3 mg/l | 0
nonhomogenous fluid in abdominal cavity | 0
fine needle aspiration from pelvis minor | 0
reddish cloudy fluid obtained | 0
diagnosis of acute peritonitis | 0
diagnostic laparoscopy | 0
peritoneal washing and drainage | 0
intraoperative esofagogastroduodenoscopy | 0
gastric-band-related defect in stomach wall | 0
purulent exudate | 0
gastric band not removed | 0
no radical surgical interventions | 0
antimicrobial therapy with Meropenem | 0
Streptococcus pyogenes (group A beta-hemolytic streptococcus) | 24
CRP level decreased | 168
discharged on 14th postoperative day | 168
readmitted to hospital at 37 weeks' gestation | 840
no complaints on admission | 840
weight 7 kg more than previous hospitalization | 840
decision not to prolong pregnancy | 840
uneventful caesarean section | 840
male neonate weighing 3060 g | 840
Apgar scores 9 at 1 min | 840
Apgar scores 10 at 5 min | 840
observed in ICU for 24 h | 840
postoperative period uneventful | 864
discharged | 864