44 years old | 0
male | 0
admitted to the hospital | 0
complaints of right lower-extremity pain | -8
progressive right lower-extremity pain | -8
untreated atrial fibrillation | 0
ulcerative colitis | 0
ongoing treatment with mesalamine | 0
agitated | 0
unable to get comfortable | 0
severe right lower-extremity pain | 0
diaphoretic | 0
tachycardic | 0
hypertensive | 0
afebrile | 0
edematous right lower extremity | 0
pulseless right lower extremity | 0
insensate right lower extremity | 0
no crepitus | 0
concern for deep vein thrombosis | 0
workup for pulmonary embolism | 0
stat computed tomography pulmonary angiogram | 0
right lower-extremity crepitus | 1
chest CT extended | 1
general surgery consulted | 1
large amount of intramuscular and intrafascial air | 1
colonic wall thickening | 1
contained perforation | 1
decision to urgently take the patient to the operating room | 1
cardiac arrest | 2
resuscitated | 2
stabilized | 2
exploratory laparotomy | 2
fasciotomy | 2
possible amputation or disarticulation | 2
subtotal colectomy | 3
pneumatosis | 3
signs of contained colonic perforation | 3
induration | 3
omental stranding | 3
hemorrhagic retroperitoneum | 3
friable retroperitoneum | 3
urology evaluation | 3
scrotum and perineum appeared healthy | 3
repositioned for orthopedic surgery | 3
numerous blisters on right lower extremity | 3
incision over proximal right thigh | 3
audible hissing of gas | 3
visible gas bubbles | 3
foul-smelling odor | 3
necrotic muscle | 3
no notable active bleeding | 3
hip disarticulated | 3
extremity placed in pathology specimen tray | 3
cultures of devitalized tissues sent | 3
necrotic muscle debulked | 3
transferred to intensive care unit | 4
multiple vasopressors | 4
multiorgan failure | 6
succumbed to multiorgan failure | 6
tissue cultures demonstrated Clostridium septicum | 6
pathology of colectomy specimen demonstrated low-grade mucinous carcinoma | 6
metastatic deposits in omentum | 6
gas gangrene | 6
necrotizing soft-tissue infection | 6
immunosuppression | 0
diabetes | 0
cancer | 0
vascular disease | 0
trauma | 0
surgery | 0
hyperbaric oxygen | 0
intravenous antibiotics | 2
debride devitalized tissue | 2
disarticulation | 3
augmentation with hyperbaric oxygen | 0
in vitro data | 0
bactericidal effects of hyperoxia | 0
emergency department room visits | 0
imaging | 0
clinical symptoms of gas gangrene | 0
radiologist | 0
diagnosis | 1
high index of suspicion | 0
early diagnosis | 0
treatment | 2
survival | 0