18 years old | 0
male | 0
chronic eczema | -720
previous alcohol abuse | -720
gout | -720
hypothyroidism | -720
presented to the emergency department | 0
worsening eruption | 0
intermittent diarrhea | 0
cutaneous eruption began | -240
desquamation of the hands | -240
desquamation of the feet | -240
perioral and perineal skin with associated pain and swelling | -240
hair loss | -240
increasing weakness | -480
fatigue | -480
70 pounds of unintentional weight loss | -480
1 to 2 glasses of wine a day | -720
smoking | -720
no significant family history | 0
not on any medications | 0
erythematous desquamative patches | 0
erosions | 0
crusted lesions | 0
diffuse nonscarring  | 0
alopecia of the scalp | 0
scaling patches on the vermillion lips | 0
methicillin-resistant Staphylococcus aureus | 0
Escherichia coli sepsis | 0
pneumonia | 0
admitted to the intensive care unit | 0
ventilator respiratory support | 0
systemic antibiotics | 0
laboratory and imaging studies | 0
ruling out necrolytic acral erythema | 0
ruling out pellagra | 0
ruling out biotin deficiency | 0
zinc levels were low | 0
antitransglutaminase and antiendomysium antibodies were positive | 0
diagnosed with celiac disease | 0
diagnosed with zinc deficiency | 0
treated with a gluten-free diet | 0
treated with zinc sulfate | 0
resolution of gastrointestinal and cutaneous symptoms | 24
acquired acrodermatitis enteropathica | -720
autosomal recessive metabolic disorder | -720
zinc transporter protein loss of function mutation | -720
SLC39A4 gene on chromosome 9 | -720
periorificial and acral dermatitis | -720
alopecia | -720
diarrhea | -720
epidermal necrosis on histology | -720
anorexia nervosa | -720
alcoholism | -720
intestinal malabsorption | -720
diets high in mineral binding phytate | -720
low zinc intake | -720
proton-pump inhibitors | -720
decreased consumption of meat and fish | -720
diets abundant in phytate-rich foods | -720
cellular and systemic zinc levels are tightly regulated | -720
anatomic sites involved in zinc homeostasis | -720
small intestine is the central avenue for homeostasis | -720
gastrointestinal pathologies decrease the absorption of zinc | -720
celiac disease | -720
inability to tolerate gliadin | -720
alcohol-soluble fraction of gluten | -720
immunologically mediated inflammatory response | -720
damage of the intestinal mucosa | -720
comorbid malabsorption | -720
diarrhea | -720
abdominal cramps | -720
flatulence | -720
weight loss | -720
growth delay in children | -720
fatigue | -720
positive immunoglobulin A antitissue transglutaminase | 0
positive antiendomysium antibodies | 0
small bowel biopsies | 0
focal villi blunting | 0
Brunner's gland hyperplasia | 0
zinc deficiency most prevalent among a comprehensive list of vitamins and minerals | 0
zinc replacement therapy | 0
adopting a gluten-free diet | 0
resolution of gastrointestinal and cutaneous symptoms | 24
acquired acrodermatitis enteropathica | -720
zinc deficiency compromises gastrointestinal epithelial barrier function | -720
pathologic conditions such as celiac disease | -720
gastrointestinal cancer | -720
inflammatory bowel disease | -720
malabsorption | -720
food allergies | -720
zinc replacement, in addition to adopting a GFD | 0
complete resolution within 4 weeks | 24