55 years old | 0
male | 0
admitted to the hospital | 0
ureteral double J stent removal | 0
left ureteric calculus | -720
endoscopic treatment | -720
compensated chronic renal failure | -8760
daily diuresis of 2500 cc volume | -8760
ureteroscopic intervention | -720
normal liver function tests | 0
hemoglobin 7.7 gr/dL | 0
hematocrit 24% | 0
WBC count 6000/uL | 0
platelet count 250,000/uL | 0
normal PT | 0
normal aPTT | 0
bilateral reduced kidney sizes | 0
increased parenchymal echogenicity | 0
ESRD | 0
creatinin clearance 7.9 mL/min | 0
protein level 2364 mg/day | 0
hemodialysis initiation | 0
ureteric catheter removal | 48
cystoscopy under sedation | 48
operation duration 10 minutes | 48
abdominal pain | 48
left upper abdominal quadrant pain | 48
abdominal distension | 48
widespread tenderness | 48
rebound positivity | 48
defense positivity | 48
body temperature 36.5°C | 48
pulse rate 105/min | 48
respiratory rate 20/min | 48
blood pressure 85/50 mm Hg | 48
urea 119 mg/dL | 48
creatinin 4.2 mg/dL | 48
sodium 140 mmol/L | 48
potassium 4.16 mmol/L | 48
hemoglobin 6.7 gr/dL | 48
hematocrit 19.9% | 48
WBC count 8000/uL | 48
platelet count 57,000/uL | 48
PT 21.7 s | 48
aPTT 110 s | 48
INR 1.91 | 48
retroperitoneal hematoma | 48
emergency exploratory operation | 48
free hemorrhagic fluid in abdomen | 48
splenic capsular laceration | 48
splenectomy | 48
fresh whole blood transfusion | 48
fresh frozen plasma transfusion | 48
thrombocyte suspension transfusion | 48
persistent thrombocytopenia | 48
high INR | 48
uremic coagulopathy diagnosis | 48
platelet transfusion | 48
fresh frozen plasma replacement | 48
stabilized blood parameters | 72
pneumococcal vaccine | 72
Hib vaccine | 72
meningococcal vaccine | 72
respiratory distress | 240
high fever | 240
pulmonary thromboembolism suspected | 240
pulmonary CT angiography | 240
sputum culture positivity for Acinetobacter | 240
blood culture positivity for Acinetobacter | 240
intravenous colimycin therapy | 240
transfer to ICU | 240
persistent high fever | 240
deteriorating respiratory distress | 240
progressive hypotension | 240
oxygen therapy need | 240
sepsis with multiorgan failure | 600
death | 600
