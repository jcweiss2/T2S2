patient underwent DALK in the left eye with big bubble technique | 0
whitish infiltrates along the graft-host junction almost 180° with severe anterior chamber reaction | 24
graft was removed and replaced by another stromal graft | 24
topical vancomycin and ceftazidime were started | 27
Gram-stain showed presence of Gram-negative Bacilli | 30
infiltrates along the entire graft host junction and hypopyon | 48
topical antibiotics were increased to half hourly | 48
report of the corneal scrapings and corneal button revealed Klebsiella pneumoniae | 72
imipenem drops was started | 72
infiltration extended toward center of graft and hypopyon persisted | 120
therapeutic penetrating keratoplasty was carried out | 120
infiltrates were observed also in host DM | 120
graft was clear without infiltrates or hypopyon | 144
gatifloxacin drops was added | 144
prednisolone drops was added | 168
unaided vision was 6/60 improving to 6/18 with pin hole | 1008
graft was clear, anterior segment was quiet with normal intraocular pressure and eradication of the pathogen | 1008
donor cornea was recovered | -6
donor cornea was preserved in McCarey Kaufman media | -72
donor cornea was transplanted | 0 
air microbiology of operation theatre was taken | 48
swabs were taken from microscope, operating tables and chairs | 48
autoclaved surgical instruments and gowns were checked | 48 
fellow donor cornea was transplanted to another recipient | 0 
patient was declared healthy | 0 
donor was declared dead | -6 
donor hospital acquired contamination of the corneal tissue | -72